//Alpha = 0. Cost: LUTs = 2859. DSPs = 144.  

`timescale 1ns / 1ps
    module mult(
        input[122:0] IN1,
        input[122:0] IN2,
        output[245:0] OUTPUT
    );
wire [16:0] slice_122;
wire [61:0] mul_55;
wire [15:0] slice_110;
wire [64:0] concat_43;
wire [31:0] mul_98;
wire [31:0] mul_31;
wire [121:0] concat_86;
wire [94:0] addW_141;
wire [16:0] addW_74;
wire [30:0] slice_7;
wire [91:0] concat_62;
wire [16:0] addW_105;
wire [33:0] mul_38;
wire [31:0] slice_93;
wire [15:0] slice_26;
wire [245:0] concat_148;
wire [64:0] concat_81;
wire [30:0] slice_14;
wire [49:0] addW_136;
wire [15:0] slice_69;
wire [15:0] slice_124;
wire [29:0] slice_57;
wire [30:0] slice_112;
wire [62:0] subW_45;
wire [15:0] slice_100;
wire [47:0] concat_33;
wire [60:0] slice_88;
wire [125:0] concat_143;
wire [33:0] mul_76;
wire [61:0] slice_9;
wire [17:0] addW_131;
wire [31:0] addW_64;
wire [32:0] addW_119;
wire [30:0] slice_52;
wire [32:0] subW_107;
wire [32:0] subW_40;
wire [62:0] addW_95;
wire [61:0] subW_83;
wire [61:0] mul_16;
wire [65:0] concat_138;
wire [31:0] mul_71;
wire [31:0] mul_126;
wire [59:0] mul_59;
wire [61:0] mul_114;
wire [30:0] slice_47;
wire [15:0] slice_102;
wire [31:0] addW_23;
wire [123:0] subW_145;
wire [32:0] subW_78;
wire [61:0] mul_11;
wire [35:0] mul_133;
wire [31:0] addW_66;
wire [32:0] addW_121;
wire [30:0] slice_54;
wire [48:0] addW_109;
wire [15:0] slice_42;
wire [15:0] slice_97;
wire [15:0] slice_30;
wire [29:0] slice_85;
wire [92:0] concat_18;
wire [63:0] subW_140;
wire [47:0] concat_73;
wire [61:0] slice_6;
wire [49:0] concat_128;
wire [29:0] slice_61;
wire [95:0] concat_116;
wire [16:0] addW_104;
wire [16:0] addW_37;
wire [62:0] addW_92;
wire [31:0] addW_25;
wire [60:0] slice_147;
wire [15:0] slice_80;
wire [33:0] subW_135;
wire [31:0] mul_68;
wire [33:0] mul_123;
wire [64:0] concat_111;
wire [62:0] subW_44;
wire [15:0] slice_99;
wire [15:0] slice_32;
wire [30:0] slice_142;
wire [16:0] addW_75;
wire [60:0] slice_51;
wire [33:0] mul_106;
wire [32:0] subW_39;
wire [15:0] slice_94;
wire [31:0] mul_27;
wire [61:0] subW_82;
wire [30:0] slice_15;
wire [15:0] slice_137;
wire [15:0] slice_70;
wire [15:0] slice_125;
wire [29:0] slice_58;
wire [30:0] slice_113;
wire [93:0] addW_46;
wire [31:0] mul_101;
wire [185:0] concat_89;
wire [123:0] subW_144;
wire [32:0] subW_77;
wire [30:0] slice_10;
wire [17:0] addW_132;
wire [15:0] slice_65;
wire [16:0] slice_120;
wire [60:0] slice_53;
wire [32:0] subW_108;
wire [48:0] addW_41;
wire [31:0] slice_96;
wire [15:0] slice_29;
wire [91:0] addW_84;
wire [30:0] slice_17;
wire [63:0] subW_139;
wire [15:0] slice_72;
wire [15:0] slice_127;
wire [30:0] slice_115;
wire [124:0] concat_48;
wire [47:0] concat_103;
wire [16:0] addW_36;
wire [15:0] slice_24;
wire [184:0] addW_146;
wire [48:0] addW_79;
wire [33:0] subW_134;
wire [15:0] slice_67;
assign slice_122 = addW_121[32:16];
assign mul_55 = slice_52 * slice_54;
assign slice_110 = mul_101[15:0];
assign concat_43 = {addW_41,slice_42};
assign mul_98 = slice_94 * slice_97;
assign mul_31 = slice_29 * slice_30;
assign concat_86 = {addW_84,slice_85};
assign addW_141 = concat_116 + subW_140;
assign addW_74 = slice_69 + slice_65;
assign slice_7 = slice_6[61:31];
assign concat_62 = {mul_55,slice_61};
assign addW_105 = slice_100 + slice_97;
assign mul_38 = addW_36 * addW_37;
assign slice_93 = addW_92[62:31];
assign slice_26 = addW_25[31:16];
assign concat_148 = {addW_146,slice_147};
assign concat_81 = {addW_79,slice_80};
assign slice_14 = slice_6[30:0];
assign addW_136 = concat_128 + subW_135;
assign slice_69 = addW_64[15:0];
assign slice_124 = addW_119[15:0];
assign slice_57 = slice_51[29:0];
assign slice_112 = addW_92[30:0];
assign subW_45 = subW_44 - mul_16;
assign slice_100 = slice_96[15:0];
assign concat_33 = {mul_27,slice_32};
assign slice_88 = concat_86[121:61];
assign concat_143 = {addW_141,slice_142};
assign mul_76 = addW_74 * addW_75;
assign slice_9 = IN2[122:61];
assign addW_131 = slice_124 + slice_120;
assign addW_64 = slice_57 + slice_52;
assign addW_119 = slice_112 + slice_93;
assign slice_52 = slice_51[60:30];
assign subW_107 = mul_106 - mul_98;
assign subW_40 = subW_39 - mul_31;
assign addW_95 = slice_53 + slice_9;
assign subW_83 = subW_82 - mul_59;
assign mul_16 = slice_14 * slice_15;
assign concat_138 = {addW_136,slice_137};
assign mul_71 = slice_69 * slice_70;
assign mul_126 = slice_124 * slice_125;
assign mul_59 = slice_57 * slice_58;
assign mul_114 = slice_112 * slice_113;
assign slice_47 = mul_16[30:0];
assign slice_102 = mul_101[31:16];
assign addW_23 = slice_14 + slice_7;
assign subW_145 = subW_144 - concat_86;
assign subW_78 = subW_77 - mul_71;
assign mul_11 = slice_7 * slice_10;
assign mul_133 = addW_131 * addW_132;
assign addW_66 = slice_58 + slice_54;
assign addW_121 = slice_113 + slice_96;
assign slice_54 = slice_53[60:30];
assign addW_109 = concat_103 + subW_108;
assign slice_42 = mul_31[15:0];
assign slice_97 = slice_96[31:16];
assign slice_30 = addW_25[15:0];
assign slice_85 = mul_59[29:0];
assign concat_18 = {mul_11,slice_17};
assign subW_140 = subW_139 - mul_114;
assign concat_73 = {mul_68,slice_72};
assign slice_6 = IN1[122:61];
assign concat_128 = {mul_123,slice_127};
assign slice_61 = mul_59[59:30];
assign concat_116 = {concat_111,slice_115};
assign addW_104 = slice_99 + slice_94;
assign addW_37 = slice_30 + slice_26;
assign addW_92 = slice_51 + slice_6;
assign addW_25 = slice_15 + slice_10;
assign slice_147 = concat_86[60:0];
assign slice_80 = mul_71[15:0];
assign subW_135 = subW_134 - mul_126;
assign mul_68 = slice_65 * slice_67;
assign mul_123 = slice_120 * slice_122;
assign concat_111 = {addW_109,slice_110};
assign subW_44 = concat_43 - mul_11;
assign slice_99 = slice_93[15:0];
assign slice_32 = mul_31[31:16];
assign slice_142 = mul_114[30:0];
assign addW_75 = slice_70 + slice_67;
assign slice_51 = IN1[60:0];
assign mul_106 = addW_104 * addW_105;
assign subW_39 = mul_38 - mul_27;
assign slice_94 = slice_93[31:16];
assign mul_27 = slice_24 * slice_26;
assign subW_82 = concat_81 - mul_55;
assign slice_15 = slice_9[30:0];
assign slice_137 = mul_126[15:0];
assign slice_70 = addW_66[15:0];
assign slice_125 = addW_121[15:0];
assign slice_58 = slice_53[29:0];
assign slice_113 = addW_95[30:0];
assign addW_46 = concat_18 + subW_45;
assign mul_101 = slice_99 * slice_100;
assign concat_89 = {concat_48,slice_88};
assign subW_144 = concat_143 - concat_48;
assign subW_77 = mul_76 - mul_68;
assign slice_10 = slice_9[61:31];
assign addW_132 = slice_125 + slice_122;
assign slice_65 = addW_64[31:16];
assign slice_120 = addW_119[32:16];
assign slice_53 = IN2[60:0];
assign subW_108 = subW_107 - mul_101;
assign addW_41 = concat_33 + subW_40;
assign slice_96 = addW_95[62:31];
assign slice_29 = addW_23[15:0];
assign addW_84 = concat_62 + subW_83;
assign slice_17 = mul_16[61:31];
assign subW_139 = concat_138 - concat_111;
assign slice_72 = mul_71[31:16];
assign slice_127 = mul_126[31:16];
assign slice_115 = mul_114[61:31];
assign concat_48 = {addW_46,slice_47};
assign concat_103 = {mul_98,slice_102};
assign addW_36 = slice_29 + slice_24;
assign slice_24 = addW_23[31:16];
assign addW_146 = concat_89 + subW_145;
assign addW_79 = concat_73 + subW_78;
assign subW_134 = mul_133 - mul_123;
assign slice_67 = addW_66[31:16];
assign OUTPUT = concat_148;
    endmodule