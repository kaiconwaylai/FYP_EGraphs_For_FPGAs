//Alpha = 0.003. Cost: LUTs = 738. DSPs = 1. 

`timescale 1ns / 1ps
    module mult(
        input[31:0] IN1,
        input[31:0] IN2,
        output[63:0] OUTPUT
    );
wire [8:0] slice_61;
wire [9:0] mul_55;
wire [4:0] slice_49;
wire [19:0] addW_43;
wire [66:0] concat_98;
wire [8:0] slice_92;
wire [6:0] slice_25;
wire [15:0] lsl_86;
wire [20:0] concat_19;
wire [8:0] mulnw_80;
wire [10:0] add_74;
wire [3:0] slice_68;
wire [8:0] slice_62;
wire [11:0] addW_56;
wire [9:0] mul_50;
wire [9:0] slice_44;
wire [17:0] slice_32;
wire [40:0] concat_93;
wire [29:0] concat_26;
wire [9:0] mul_87;
wire [18:0] lsl_81;
wire [15:0] lsl_75;
wire [6:0] slice_8;
wire [8:0] mulnw_69;
wire [17:0] mul_63;
wire [16:0] addW_57;
wire [4:0] slice_51;
wire [4:0] slice_45;
wire [19:0] addW_39;
wire [47:0] concat_33;
wire [41:0] subW_94;
wire [16:0] add_88;
wire [13:0] mul_21;
wire [4:0] slice_82;
wire [6:0] slice_15;
wire [9:0] mul_76;
wire [18:0] lsl_70;
wire [8:0] slice_64;
wire [4:0] slice_58;
wire [14:0] concat_52;
wire [9:0] mul_46;
wire [42:0] subW_95;
wire [17:0] slice_28;
wire [19:0] add_89;
wire [13:0] mul_22;
wire [9:0] mulnw_83;
wire [6:0] slice_16;
wire [16:0] add_77;
wire [13:0] slice_10;
wire [8:0] mulnw_71;
wire [30:0] concat_65;
wire [21:0] concat_59;
wire [9:0] slice_41;
wire [48:0] addW_96;
wire [17:0] slice_29;
wire [20:0] addW_90;
wire [15:0] addW_23;
wire [8:0] mulnw_84;
wire [13:0] mul_17;
wire [19:0] add_78;
wire [6:0] slice_11;
wire [4:0] slice_72;
wire [9:0] mul_54;
wire [4:0] slice_48;
wire [4:0] slice_42;
wire [17:0] slice_97;
wire [35:0] mul_30;
wire [31:0] addW_91;
wire [22:0] addW_24;
wire [10:0] add_85;
wire [6:0] slice_18;
wire [3:0] slice_79;
wire [13:0] mul_12;
wire [9:0] mulnw_73;
wire [13:0] slice_6;
assign slice_61 = addW_39[8:0];
assign mul_55 = slice_48 * slice_45;
assign slice_49 = slice_44[4:0];
assign addW_43 = slice_29 + slice_10;
assign concat_98 = {addW_96,slice_97};
assign slice_92 = mul_63[8:0];
assign slice_25 = mul_17[6:0];
assign lsl_86 = add_85 << 5;
assign concat_19 = {mul_12,slice_18};
assign mulnw_80 = slice_79 * slice_45;
assign add_74 = mulnw_71 + mulnw_73;
assign slice_68 = slice_62[8:5];
assign slice_62 = addW_43[8:0];
assign addW_56 = mul_54 + mul_55;
assign mul_50 = slice_48 * slice_49;
assign slice_44 = addW_43[18:9];
assign slice_32 = mul_30[35:18];
assign concat_93 = {addW_91,slice_92};
assign concat_26 = {addW_24,slice_25};
assign mul_87 = slice_82 * slice_49;
assign lsl_81 = mulnw_80 << 10;
assign lsl_75 = add_74 << 5;
assign slice_8 = slice_6[13:7];
assign mulnw_69 = slice_42 * slice_68;
assign mul_63 = slice_61 * slice_62;
assign addW_57 = concat_52 + addW_56;
assign slice_51 = mul_50[9:5];
assign slice_45 = slice_44[9:5];
assign addW_39 = slice_28 + slice_6;
assign concat_33 = {concat_26,slice_32};
assign subW_94 = concat_93 - concat_26;
assign add_88 = lsl_86 + mul_87;
assign mul_21 = slice_8 * slice_16;
assign slice_82 = slice_61[4:0];
assign slice_15 = slice_6[6:0];
assign mul_76 = slice_48 * slice_72;
assign lsl_70 = mulnw_69 << 10;
assign slice_64 = mul_63[17:9];
assign slice_58 = mul_50[4:0];
assign concat_52 = {mul_46,slice_51};
assign mul_46 = slice_42 * slice_45;
assign subW_95 = subW_94 - mul_30;
assign slice_28 = IN1[17:0];
assign add_89 = lsl_81 + add_88;
assign mul_22 = slice_15 * slice_11;
assign mulnw_83 = slice_82 * slice_45;
assign slice_16 = slice_10[6:0];
assign add_77 = lsl_75 + mul_76;
assign slice_10 = IN2[31:18];
assign mulnw_71 = slice_48 * slice_68;
assign concat_65 = {concat_59,slice_64};
assign concat_59 = {addW_57,slice_58};
assign slice_41 = addW_39[18:9];
assign addW_96 = concat_33 + subW_95;
assign slice_29 = IN2[17:0];
assign addW_90 = add_78 + add_89;
assign addW_23 = mul_21 + mul_22;
assign mulnw_84 = slice_79 * slice_49;
assign mul_17 = slice_15 * slice_16;
assign add_78 = lsl_70 + add_77;
assign slice_11 = slice_10[13:7];
assign slice_72 = slice_62[4:0];
assign mul_54 = slice_42 * slice_49;
assign slice_48 = slice_41[4:0];
assign slice_42 = slice_41[9:5];
assign slice_97 = mul_30[17:0];
assign mul_30 = slice_28 * slice_29;
assign addW_91 = concat_65 + addW_90;
assign addW_24 = concat_19 + addW_23;
assign add_85 = mulnw_83 + mulnw_84;
assign slice_18 = mul_17[13:7];
assign slice_79 = slice_61[8:5];
assign mul_12 = slice_8 * slice_11;
assign mulnw_73 = slice_42 * slice_72;
assign slice_6 = IN1[31:18];
assign OUTPUT = concat_98;
    endmodule