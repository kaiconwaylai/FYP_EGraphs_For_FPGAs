//Alpha = 0.007. Cost: LUTs = 0. DSPs = 18.  

`timescale 1ns / 1ps
    module mult(
        input[126:0] IN1,
        input[126:0] IN2,
        output[253:0] OUTPUT
    );
wire [49:0] concat_189;
wire [7:0] slice_55;
wire [30:0] lsl_110;
wire [50:0] addW_165;
wire [15:0] slice_31;
wire [31:0] slice_220;
wire [31:0] mul_86;
wire [32:0] lsl_141;
wire [31:0] slice_7;
wire [7:0] slice_196;
wire [26:0] add_62;
wire [15:0] mul_117;
wire [126:0] concat_172;
wire [7:0] slice_38;
wire [34:0] addW_227;
wire [46:0] concat_93;
wire [15:0] mul_148;
wire [31:0] slice_14;
wire [7:0] slice_203;
wire [68:0] subW_69;
wire [32:0] slice_179;
wire [16:0] mulnw_45;
wire [132:0] subW_234;
wire [7:0] slice_100;
wire [7:0] slice_155;
wire [15:0] mulnw_210;
wire [31:0] slice_76;
wire [16:0] slice_131;
wire [15:0] slice_186;
wire [8:0] slice_52;
wire [6:0] slice_107;
wire [26:0] add_162;
wire [33:0] mul_28;
wire [50:0] addW_217;
wire [15:0] slice_83;
wire [8:0] slice_138;
wire [32:0] lsl_193;
wire [17:0] add_59;
wire [14:0] mulnw_114;
wire [68:0] subW_169;
wire [98:0] concat_224;
wire [29:0] mul_90;
wire [16:0] mulnw_145;
wire [63:0] mul_11;
wire [15:0] mul_200;
wire [15:0] slice_66;
wire [47:0] addW_121;
wire [7:0] slice_42;
wire [99:0] addW_231;
wire [30:0] lsl_97;
wire [8:0] slice_152;
wire [95:0] concat_18;
wire [7:0] slice_207;
wire [33:0] addW_128;
wire [16:0] slice_183;
wire [26:0] add_49;
wire [256:0] concat_238;
wire [15:0] mul_104;
wire [17:0] add_159;
wire [16:0] slice_25;
wire [26:0] add_214;
wire [31:0] mul_135;
wire [8:0] slice_190;
wire [16:0] mulnw_56;
wire [7:0] slice_111;
wire [15:0] slice_166;
wire [31:0] mul_32;
wire [31:0] slice_221;
wire [7:0] slice_142;
wire [16:0] mulnw_197;
wire [33:0] add_63;
wire [25:0] add_118;
wire [16:0] mulnw_39;
wire [69:0] mul_228;
wire [7:0] slice_94;
wire [26:0] add_149;
wire [31:0] slice_15;
wire [8:0] slice_204;
wire [97:0] addW_70;
wire [30:0] slice_125;
wire [16:0] slice_180;
wire [17:0] add_46;
wire [133:0] subW_235;
wire [15:0] mulnw_101;
wire [16:0] mulnw_156;
wire [17:0] add_211;
wire [62:0] slice_77;
wire [33:0] mul_132;
wire [31:0] mul_187;
wire [16:0] mulnw_53;
wire [7:0] slice_108;
wire [33:0] add_163;
wire [15:0] slice_218;
wire [30:0] slice_84;
wire [7:0] slice_139;
wire [7:0] slice_194;
wire [25:0] lsl_60;
wire [16:0] add_115;
wire [95:0] addW_170;
wire [17:0] add_146;
wire [26:0] add_201;
wire [66:0] concat_67;
wire [14:0] slice_122;
wire [15:0] mulnw_43;
wire [31:0] slice_232;
wire [7:0] slice_98;
wire [16:0] mulnw_153;
wire [16:0] mulnw_208;
wire [16:0] slice_129;
wire [33:0] mul_184;
wire [33:0] add_50;
wire [25:0] add_105;
wire [25:0] lsl_160;
wire [33:0] addW_26;
wire [33:0] add_215;
wire [15:0] slice_136;
wire [7:0] slice_191;
wire [7:0] slice_57;
wire [15:0] mulnw_112;
wire [66:0] concat_167;
wire [15:0] slice_33;
wire [63:0] mul_222;
wire [14:0] slice_88;
wire [15:0] mulnw_143;
wire [63:0] slice_9;
wire [17:0] add_198;
wire [34:0] addW_64;
wire [31:0] add_119;
wire [62:0] slice_174;
wire [32:0] lsl_40;
wire [70:0] subW_229;
wire [6:0] slice_95;
wire [33:0] add_150;
wire [63:0] mul_16;
wire [16:0] mulnw_205;
wire [31:0] slice_71;
wire [94:0] concat_126;
wire [65:0] addW_181;
wire [25:0] lsl_47;
wire [193:0] addW_236;
wire [16:0] add_102;
wire [7:0] slice_157;
wire [33:0] addW_23;
wire [25:0] lsl_212;
wire [31:0] slice_78;
wire [15:0] slice_133;
wire [15:0] slice_188;
wire [32:0] lsl_54;
wire [14:0] mulnw_109;
wire [34:0] addW_164;
wire [15:0] slice_30;
wire [66:0] concat_219;
wire [15:0] slice_85;
wire [16:0] mulnw_140;
wire [63:0] slice_6;
wire [15:0] mulnw_195;
wire [15:0] mul_61;
wire [24:0] lsl_116;
wire [30:0] slice_171;
wire [8:0] slice_37;
wire [34:0] addW_226;
wire [14:0] slice_92;
wire [25:0] lsl_147;
wire [33:0] add_202;
wire [67:0] subW_68;
wire [62:0] concat_123;
wire [65:0] addW_178;
wire [7:0] slice_44;
wire [131:0] concat_233;
wire [14:0] mulnw_99;
wire [32:0] lsl_154;
wire [7:0] slice_209;
wire [62:0] slice_75;
wire [33:0] addW_130;
wire [15:0] slice_185;
wire [7:0] slice_51;
wire [31:0] add_106;
wire [15:0] mul_161;
wire [16:0] slice_27;
wire [34:0] addW_216;
wire [30:0] slice_82;
wire [49:0] concat_137;
wire [16:0] mulnw_192;
wire [15:0] mulnw_58;
wire [7:0] slice_113;
wire [67:0] subW_168;
wire [49:0] concat_34;
wire [31:0] slice_223;
wire [14:0] slice_89;
wire [7:0] slice_144;
wire [31:0] slice_10;
wire [25:0] lsl_199;
wire [50:0] addW_65;
wire [32:0] addW_120;
wire [192:0] concat_175;
wire [71:0] subW_230;
wire [14:0] mulnw_96;
wire [7:0] slice_151;
wire [31:0] slice_17;
wire [32:0] lsl_206;
wire [129:0] concat_72;
wire [32:0] slice_182;
wire [15:0] mul_48;
wire [62:0] slice_237;
wire [24:0] lsl_103;
wire [15:0] mulnw_158;
wire [15:0] mul_213;
wire [63:0] mul_79;
wire [15:0] slice_134;
assign concat_189 = {mul_184,slice_188};
assign slice_55 = slice_30[7:0];
assign lsl_110 = mulnw_109 << 16;
assign addW_165 = concat_137 + addW_164;
assign slice_31 = addW_26[15:0];
assign slice_220 = addW_178[31:0];
assign mul_86 = slice_83 * slice_85;
assign lsl_141 = mulnw_140 << 16;
assign slice_7 = slice_6[63:32];
assign slice_196 = slice_186[7:0];
assign add_62 = lsl_60 + mul_61;
assign mul_117 = slice_111 * slice_113;
assign concat_172 = {addW_170,slice_171};
assign slice_38 = slice_31[15:8];
assign addW_227 = slice_221 + slice_182;
assign concat_93 = {mul_86,slice_92};
assign mul_148 = slice_142 * slice_144;
assign slice_14 = slice_6[31:0];
assign slice_203 = slice_185[15:8];
assign subW_69 = subW_68 - mul_16;
assign slice_179 = addW_178[64:32];
assign mulnw_45 = slice_37 * slice_44;
assign subW_234 = concat_233 - concat_72;
assign slice_100 = slice_89[7:0];
assign slice_155 = slice_133[7:0];
assign mulnw_210 = slice_203 * slice_209;
assign slice_76 = slice_75[62:31];
assign slice_131 = addW_130[32:16];
assign slice_186 = slice_182[15:0];
assign slice_52 = slice_27[16:8];
assign slice_107 = slice_88[14:8];
assign add_162 = lsl_160 + mul_161;
assign mul_28 = slice_25 * slice_27;
assign addW_217 = concat_189 + addW_216;
assign slice_83 = slice_82[30:15];
assign slice_138 = slice_129[16:8];
assign lsl_193 = mulnw_192 << 16;
assign add_59 = mulnw_56 + mulnw_58;
assign mulnw_114 = slice_107 * slice_113;
assign subW_169 = subW_168 - concat_123;
assign concat_224 = {concat_219,slice_223};
assign mul_90 = slice_88 * slice_89;
assign mulnw_145 = slice_138 * slice_144;
assign mul_11 = slice_7 * slice_10;
assign mul_200 = slice_194 * slice_196;
assign slice_66 = mul_32[15:0];
assign addW_121 = concat_93 + addW_120;
assign slice_42 = slice_25[7:0];
assign addW_231 = concat_224 + subW_230;
assign lsl_97 = mulnw_96 << 16;
assign slice_152 = slice_131[16:8];
assign concat_18 = {mul_11,slice_17};
assign slice_207 = slice_185[7:0];
assign addW_128 = slice_82 + slice_76;
assign slice_183 = slice_182[32:16];
assign add_49 = lsl_47 + mul_48;
assign concat_238 = {addW_236,slice_237};
assign mul_104 = slice_98 * slice_100;
assign add_159 = mulnw_156 + mulnw_158;
assign slice_25 = addW_23[32:16];
assign add_214 = lsl_212 + mul_213;
assign mul_135 = slice_133 * slice_134;
assign slice_190 = slice_180[16:8];
assign mulnw_56 = slice_55 * slice_52;
assign slice_111 = slice_88[7:0];
assign slice_166 = mul_135[15:0];
assign mul_32 = slice_30 * slice_31;
assign slice_221 = addW_181[31:0];
assign slice_142 = slice_129[7:0];
assign mulnw_197 = slice_190 * slice_196;
assign add_63 = lsl_54 + add_62;
assign add_118 = lsl_116 + mul_117;
assign mulnw_39 = slice_37 * slice_38;
assign mul_228 = addW_226 * addW_227;
assign slice_94 = slice_83[15:8];
assign add_149 = lsl_147 + mul_148;
assign slice_15 = slice_9[31:0];
assign slice_204 = slice_183[16:8];
assign addW_70 = concat_18 + subW_69;
assign slice_125 = concat_123[61:31];
assign slice_180 = slice_179[32:16];
assign add_46 = mulnw_43 + mulnw_45;
assign subW_235 = subW_234 - concat_172;
assign mulnw_101 = slice_94 * slice_100;
assign mulnw_156 = slice_155 * slice_152;
assign add_211 = mulnw_208 + mulnw_210;
assign slice_77 = IN2[62:0];
assign mul_132 = slice_129 * slice_131;
assign mul_187 = slice_185 * slice_186;
assign mulnw_53 = slice_51 * slice_52;
assign slice_108 = slice_85[15:8];
assign add_163 = lsl_154 + add_162;
assign slice_218 = mul_187[15:0];
assign slice_84 = slice_77[30:0];
assign slice_139 = slice_134[15:8];
assign slice_194 = slice_180[7:0];
assign lsl_60 = add_59 << 8;
assign add_115 = mulnw_112 + mulnw_114;
assign addW_170 = concat_126 + subW_169;
assign add_146 = mulnw_143 + mulnw_145;
assign add_201 = lsl_199 + mul_200;
assign concat_67 = {addW_65,slice_66};
assign slice_122 = mul_90[14:0];
assign mulnw_43 = slice_42 * slice_38;
assign slice_232 = mul_222[31:0];
assign slice_98 = slice_83[7:0];
assign mulnw_153 = slice_151 * slice_152;
assign mulnw_208 = slice_207 * slice_204;
assign slice_129 = addW_128[32:16];
assign mul_184 = slice_180 * slice_183;
assign add_50 = lsl_40 + add_49;
assign add_105 = lsl_103 + mul_104;
assign lsl_160 = add_159 << 8;
assign addW_26 = slice_15 + slice_10;
assign add_215 = lsl_206 + add_214;
assign slice_136 = mul_135[31:16];
assign slice_191 = slice_186[15:8];
assign slice_57 = slice_27[7:0];
assign mulnw_112 = slice_111 * slice_108;
assign concat_167 = {addW_165,slice_166};
assign slice_33 = mul_32[31:16];
assign mul_222 = slice_220 * slice_221;
assign slice_88 = slice_82[14:0];
assign mulnw_143 = slice_142 * slice_139;
assign slice_9 = IN2[126:63];
assign add_198 = mulnw_195 + mulnw_197;
assign addW_64 = add_50 + add_63;
assign add_119 = lsl_110 + add_118;
assign slice_174 = concat_172[125:63];
assign lsl_40 = mulnw_39 << 16;
assign subW_229 = mul_228 - concat_219;
assign slice_95 = slice_89[14:8];
assign add_150 = lsl_141 + add_149;
assign mul_16 = slice_14 * slice_15;
assign mulnw_205 = slice_203 * slice_204;
assign slice_71 = mul_16[31:0];
assign concat_126 = {mul_79,slice_125};
assign addW_181 = slice_77 + slice_9;
assign lsl_47 = add_46 << 8;
assign addW_236 = concat_175 + subW_235;
assign add_102 = mulnw_99 + mulnw_101;
assign slice_157 = slice_131[7:0];
assign addW_23 = slice_14 + slice_7;
assign lsl_212 = add_211 << 8;
assign slice_78 = slice_77[62:31];
assign slice_133 = addW_128[15:0];
assign slice_188 = mul_187[31:16];
assign lsl_54 = mulnw_53 << 16;
assign mulnw_109 = slice_107 * slice_108;
assign addW_164 = add_150 + add_163;
assign slice_30 = addW_23[15:0];
assign concat_219 = {addW_217,slice_218};
assign slice_85 = slice_84[30:15];
assign mulnw_140 = slice_138 * slice_139;
assign slice_6 = IN1[126:63];
assign mulnw_195 = slice_194 * slice_191;
assign mul_61 = slice_55 * slice_57;
assign lsl_116 = add_115 << 8;
assign slice_171 = concat_123[30:0];
assign slice_37 = slice_25[16:8];
assign addW_226 = slice_220 + slice_179;
assign slice_92 = mul_90[29:15];
assign lsl_147 = add_146 << 8;
assign add_202 = lsl_193 + add_201;
assign subW_68 = concat_67 - mul_11;
assign concat_123 = {addW_121,slice_122};
assign addW_178 = slice_75 + slice_6;
assign slice_44 = slice_31[7:0];
assign concat_233 = {addW_231,slice_232};
assign mulnw_99 = slice_98 * slice_95;
assign lsl_154 = mulnw_153 << 16;
assign slice_209 = slice_183[7:0];
assign slice_75 = IN1[62:0];
assign addW_130 = slice_84 + slice_78;
assign slice_185 = slice_179[15:0];
assign slice_51 = slice_30[15:8];
assign add_106 = lsl_97 + add_105;
assign mul_161 = slice_155 * slice_157;
assign slice_27 = addW_26[32:16];
assign addW_216 = add_202 + add_215;
assign slice_82 = slice_75[30:0];
assign concat_137 = {mul_132,slice_136};
assign mulnw_192 = slice_190 * slice_191;
assign mulnw_58 = slice_51 * slice_57;
assign slice_113 = slice_85[7:0];
assign subW_168 = concat_167 - mul_79;
assign concat_34 = {mul_28,slice_33};
assign slice_223 = mul_222[63:32];
assign slice_89 = slice_84[14:0];
assign slice_144 = slice_134[7:0];
assign slice_10 = slice_9[63:32];
assign lsl_199 = add_198 << 8;
assign addW_65 = concat_34 + addW_64;
assign addW_120 = add_106 + add_119;
assign concat_175 = {concat_72,slice_174};
assign subW_230 = subW_229 - mul_222;
assign mulnw_96 = slice_94 * slice_95;
assign slice_151 = slice_133[15:8];
assign slice_17 = mul_16[63:32];
assign lsl_206 = mulnw_205 << 16;
assign concat_72 = {addW_70,slice_71};
assign slice_182 = addW_181[64:32];
assign mul_48 = slice_42 * slice_44;
assign slice_237 = concat_172[62:0];
assign lsl_103 = add_102 << 8;
assign mulnw_158 = slice_151 * slice_157;
assign mul_213 = slice_207 * slice_209;
assign mul_79 = slice_76 * slice_78;
assign slice_134 = addW_130[15:0];
assign OUTPUT = concat_238;
    endmodule