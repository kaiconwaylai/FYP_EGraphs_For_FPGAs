Alpha = 0.003. Cost: LUTs = 2321. DSPs = 3. 

`timescale 1ns / 1ps
    module mult(
        input[63:0] IN1,
        input[63:0] IN2,
        output[127:0] OUTPUT
    );
wire [16:0] slice_189;
wire [9:0] mul_55;
wire [13:0] mul_110;
wire [9:0] mulnw_165;
wire [29:0] concat_31;
wire [26:0] add_220;
wire [18:0] lsl_86;
wire [11:0] addW_141;
wire [31:0] slice_7;
wire [15:0] mul_196;
wire [16:0] addW_62;
wire [13:0] mul_117;
wire [20:0] addW_172;
wire [47:0] concat_38;
wire [15:0] mulnw_227;
wire [16:0] add_93;
wire [8:0] slice_148;
wire [31:0] slice_14;
wire [15:0] mul_203;
wire [8:0] slice_69;
wire [35:0] mul_124;
wire [17:0] slice_179;
wire [50:0] addW_234;
wire [42:0] subW_100;
wire [9:0] mulnw_155;
wire [6:0] slice_21;
wire [8:0] mulnw_76;
wire [9:0] slice_131;
wire [33:0] addW_186;
wire [131:0] concat_241;
wire [31:0] slice_107;
wire [8:0] mulnw_162;
wire [15:0] addW_28;
wire [17:0] add_217;
wire [19:0] add_83;
wire [14:0] concat_138;
wire [7:0] slice_193;
wire [9:0] mul_59;
wire [6:0] slice_114;
wire [9:0] mul_169;
wire [35:0] mul_35;
wire [32:0] lsl_224;
wire [10:0] add_90;
wire [8:0] slice_145;
wire [7:0] slice_200;
wire [8:0] slice_66;
wire [29:0] concat_121;
wire [41:0] subW_176;
wire [26:0] add_231;
wire [8:0] slice_97;
wire [18:0] lsl_152;
wire [33:0] concat_207;
wire [3:0] slice_73;
wire [9:0] slice_128;
wire [9:0] slice_49;
wire [68:0] subW_238;
wire [31:0] slice_104;
wire [16:0] add_159;
wire [7:0] slice_214;
wire [15:0] lsl_80;
wire [4:0] slice_135;
wire [33:0] mul_190;
wire [4:0] slice_56;
wire [6:0] slice_111;
wire [8:0] mulnw_166;
wire [33:0] add_221;
wire [4:0] slice_87;
wire [16:0] addW_142;
wire [7:0] slice_197;
wire [4:0] slice_63;
wire [15:0] addW_118;
wire [31:0] addW_173;
wire [17:0] add_228;
wire [19:0] add_94;
wire [30:0] concat_149;
wire [13:0] slice_15;
wire [17:0] addW_204;
wire [30:0] concat_70;
wire [17:0] slice_125;
wire [66:0] concat_180;
wire [9:0] slice_46;
wire [15:0] slice_235;
wire [48:0] addW_101;
wire [10:0] add_156;
wire [13:0] mul_22;
wire [8:0] slice_211;
wire [4:0] slice_77;
wire [4:0] slice_132;
wire [16:0] slice_187;
wire [4:0] slice_53;
wire [13:0] slice_108;
wire [18:0] lsl_163;
wire [22:0] addW_29;
wire [25:0] lsl_218;
wire [3:0] slice_84;
wire [9:0] mul_139;
wire [15:0] slice_194;
wire [9:0] mul_60;
wire [20:0] concat_115;
wire [16:0] add_170;
wire [16:0] mulnw_225;
wire [15:0] lsl_91;
wire [8:0] slice_146;
wire [6:0] slice_12;
wire [23:0] concat_201;
wire [8:0] slice_67;
wire [17:0] slice_122;
wire [42:0] subW_177;
wire [33:0] add_232;
wire [40:0] concat_98;
wire [8:0] mulnw_153;
wire [15:0] slice_208;
wire [8:0] mulnw_74;
wire [4:0] slice_129;
wire [4:0] slice_50;
wire [99:0] addW_239;
wire [13:0] slice_105;
wire [19:0] add_160;
wire [13:0] mul_26;
wire [15:0] mulnw_215;
wire [9:0] mul_81;
wire [9:0] mul_136;
wire [14:0] concat_57;
wire [6:0] slice_112;
wire [10:0] add_167;
wire [17:0] slice_33;
wire [8:0] slice_222;
wire [9:0] mulnw_88;
wire [4:0] slice_143;
wire [7:0] slice_198;
wire [21:0] concat_64;
wire [22:0] addW_119;
wire [8:0] slice_174;
wire [25:0] lsl_229;
wire [20:0] addW_95;
wire [3:0] slice_150;
wire [6:0] slice_16;
wire [25:0] addW_205;
wire [47:0] concat_126;
wire [31:0] slice_181;
wire [4:0] slice_47;
wire [66:0] concat_236;
wire [17:0] slice_102;
wire [15:0] lsl_157;
wire [6:0] slice_23;
wire [16:0] mulnw_212;
wire [9:0] mulnw_78;
wire [9:0] mul_133;
wire [33:0] addW_188;
wire [4:0] slice_54;
wire [6:0] slice_109;
wire [4:0] slice_164;
wire [6:0] slice_30;
wire [15:0] mul_219;
wire [8:0] mulnw_85;
wire [9:0] mul_140;
wire [7:0] slice_195;
wire [11:0] addW_61;
wire [13:0] mul_116;
wire [19:0] add_171;
wire [17:0] slice_37;
wire [7:0] slice_226;
wire [9:0] mul_92;
wire [17:0] mul_147;
wire [15:0] mul_202;
wire [17:0] mul_68;
wire [17:0] slice_123;
wire [48:0] addW_178;
wire [19:0] addW_44;
wire [34:0] addW_233;
wire [41:0] subW_99;
wire [4:0] slice_154;
wire [6:0] slice_20;
wire [49:0] concat_209;
wire [18:0] lsl_75;
wire [19:0] addW_130;
wire [9:0] mul_51;
wire [31:0] slice_240;
wire [6:0] slice_106;
wire [3:0] slice_161;
wire [13:0] mul_27;
wire [16:0] mulnw_216;
wire [16:0] add_82;
wire [4:0] slice_137;
wire [15:0] slice_192;
wire [13:0] mul_113;
wire [15:0] lsl_168;
wire [17:0] slice_34;
wire [16:0] mulnw_223;
wire [8:0] mulnw_89;
wire [21:0] concat_144;
wire [13:0] slice_10;
wire [15:0] mul_199;
wire [6:0] slice_120;
wire [40:0] concat_175;
wire [15:0] mul_230;
wire [31:0] addW_96;
wire [8:0] mulnw_151;
wire [13:0] mul_17;
wire [7:0] slice_206;
wire [19:0] addW_127;
wire [98:0] concat_182;
wire [19:0] addW_48;
wire [67:0] subW_237;
wire [66:0] concat_103;
wire [9:0] mul_158;
wire [20:0] concat_24;
wire [32:0] lsl_213;
wire [10:0] add_79;
wire [4:0] slice_134;
assign slice_189 = addW_188[32:16];
assign mul_55 = slice_53 * slice_54;
assign mul_110 = slice_106 * slice_109;
assign mulnw_165 = slice_164 * slice_132;
assign concat_31 = {addW_29,slice_30};
assign add_220 = lsl_218 + mul_219;
assign lsl_86 = mulnw_85 << 10;
assign addW_141 = mul_139 + mul_140;
assign slice_7 = IN1[63:32];
assign mul_196 = slice_193 * slice_195;
assign addW_62 = concat_57 + addW_61;
assign mul_117 = slice_111 * slice_109;
assign addW_172 = add_160 + add_171;
assign concat_38 = {concat_31,slice_37};
assign mulnw_227 = slice_193 * slice_226;
assign add_93 = lsl_91 + mul_92;
assign slice_148 = mul_147[17:9];
assign slice_14 = IN2[63:32];
assign mul_203 = slice_197 * slice_195;
assign slice_69 = mul_68[17:9];
assign mul_124 = slice_122 * slice_123;
assign slice_179 = mul_124[17:0];
assign addW_234 = concat_209 + addW_233;
assign subW_100 = subW_99 - mul_35;
assign mulnw_155 = slice_129 * slice_154;
assign slice_21 = slice_15[6:0];
assign mulnw_76 = slice_53 * slice_73;
assign slice_131 = addW_130[18:9];
assign addW_186 = slice_104 + slice_7;
assign concat_241 = {addW_239,slice_240};
assign slice_107 = IN2[31:0];
assign mulnw_162 = slice_161 * slice_132;
assign addW_28 = mul_26 + mul_27;
assign add_217 = mulnw_215 + mulnw_216;
assign add_83 = lsl_75 + add_82;
assign concat_138 = {mul_133,slice_137};
assign slice_193 = slice_192[15:8];
assign mul_59 = slice_47 * slice_54;
assign slice_114 = mul_113[13:7];
assign mul_169 = slice_164 * slice_135;
assign mul_35 = slice_33 * slice_34;
assign lsl_224 = mulnw_223 << 16;
assign add_90 = mulnw_88 + mulnw_89;
assign slice_145 = addW_127[8:0];
assign slice_200 = mul_199[15:8];
assign slice_66 = addW_44[8:0];
assign concat_121 = {addW_119,slice_120};
assign subW_176 = concat_175 - concat_121;
assign add_231 = lsl_229 + mul_230;
assign slice_97 = mul_68[8:0];
assign lsl_152 = mulnw_151 << 10;
assign concat_207 = {addW_205,slice_206};
assign slice_73 = slice_67[8:5];
assign slice_128 = addW_127[18:9];
assign slice_49 = addW_48[18:9];
assign subW_238 = subW_237 - concat_180;
assign slice_104 = IN1[31:0];
assign add_159 = lsl_157 + mul_158;
assign slice_214 = slice_187[7:0];
assign lsl_80 = add_79 << 5;
assign slice_135 = slice_131[4:0];
assign mul_190 = slice_187 * slice_189;
assign slice_56 = mul_55[9:5];
assign slice_111 = slice_105[6:0];
assign mulnw_166 = slice_161 * slice_135;
assign add_221 = lsl_213 + add_220;
assign slice_87 = slice_66[4:0];
assign addW_142 = concat_138 + addW_141;
assign slice_197 = slice_192[7:0];
assign slice_63 = mul_55[4:0];
assign addW_118 = mul_116 + mul_117;
assign addW_173 = concat_149 + addW_172;
assign add_228 = mulnw_225 + mulnw_227;
assign add_94 = lsl_86 + add_93;
assign concat_149 = {concat_144,slice_148};
assign slice_15 = slice_14[31:18];
assign addW_204 = mul_202 + mul_203;
assign concat_70 = {concat_64,slice_69};
assign slice_125 = mul_124[35:18];
assign concat_180 = {addW_178,slice_179};
assign slice_46 = addW_44[18:9];
assign slice_235 = concat_207[15:0];
assign addW_101 = concat_38 + subW_100;
assign add_156 = mulnw_153 + mulnw_155;
assign mul_22 = slice_20 * slice_21;
assign slice_211 = slice_187[16:8];
assign slice_77 = slice_67[4:0];
assign slice_132 = slice_131[9:5];
assign slice_187 = addW_186[32:16];
assign slice_53 = slice_46[4:0];
assign slice_108 = slice_107[31:18];
assign lsl_163 = mulnw_162 << 10;
assign addW_29 = concat_24 + addW_28;
assign lsl_218 = add_217 << 8;
assign slice_84 = slice_66[8:5];
assign mul_139 = slice_129 * slice_135;
assign slice_194 = addW_188[15:0];
assign mul_60 = slice_53 * slice_50;
assign concat_115 = {mul_110,slice_114};
assign add_170 = lsl_168 + mul_169;
assign mulnw_225 = slice_197 * slice_222;
assign lsl_91 = add_90 << 5;
assign slice_146 = addW_130[8:0];
assign slice_12 = slice_10[13:7];
assign concat_201 = {mul_196,slice_200};
assign slice_67 = addW_48[8:0];
assign slice_122 = slice_104[17:0];
assign subW_177 = subW_176 - mul_124;
assign add_232 = lsl_224 + add_231;
assign concat_98 = {addW_96,slice_97};
assign mulnw_153 = slice_134 * slice_150;
assign slice_208 = concat_207[31:16];
assign mulnw_74 = slice_47 * slice_73;
assign slice_129 = slice_128[9:5];
assign slice_50 = slice_49[9:5];
assign addW_239 = concat_182 + subW_238;
assign slice_105 = slice_104[31:18];
assign add_160 = lsl_152 + add_159;
assign mul_26 = slice_12 * slice_21;
assign mulnw_215 = slice_214 * slice_195;
assign mul_81 = slice_53 * slice_77;
assign mul_136 = slice_134 * slice_135;
assign concat_57 = {mul_51,slice_56};
assign slice_112 = slice_108[6:0];
assign add_167 = mulnw_165 + mulnw_166;
assign slice_33 = slice_7[17:0];
assign slice_222 = slice_189[16:8];
assign mulnw_88 = slice_87 * slice_50;
assign slice_143 = mul_136[4:0];
assign slice_198 = slice_194[7:0];
assign concat_64 = {addW_62,slice_63};
assign addW_119 = concat_115 + addW_118;
assign slice_174 = mul_147[8:0];
assign lsl_229 = add_228 << 8;
assign addW_95 = add_83 + add_94;
assign slice_150 = slice_146[8:5];
assign slice_16 = slice_15[13:7];
assign addW_205 = concat_201 + addW_204;
assign concat_126 = {concat_121,slice_125};
assign slice_181 = concat_180[63:32];
assign slice_47 = slice_46[9:5];
assign concat_236 = {addW_234,slice_235};
assign slice_102 = mul_35[17:0];
assign lsl_157 = add_156 << 5;
assign slice_23 = mul_22[13:7];
assign mulnw_212 = slice_211 * slice_195;
assign mulnw_78 = slice_47 * slice_77;
assign mul_133 = slice_129 * slice_132;
assign addW_188 = slice_107 + slice_14;
assign slice_54 = slice_49[4:0];
assign slice_109 = slice_108[13:7];
assign slice_164 = slice_145[4:0];
assign slice_30 = mul_22[6:0];
assign mul_219 = slice_214 * slice_198;
assign mulnw_85 = slice_84 * slice_50;
assign mul_140 = slice_134 * slice_132;
assign slice_195 = slice_194[15:8];
assign addW_61 = mul_59 + mul_60;
assign mul_116 = slice_106 * slice_112;
assign add_171 = lsl_163 + add_170;
assign slice_37 = mul_35[35:18];
assign slice_226 = slice_189[7:0];
assign mul_92 = slice_87 * slice_54;
assign mul_147 = slice_145 * slice_146;
assign mul_202 = slice_193 * slice_198;
assign mul_68 = slice_66 * slice_67;
assign slice_123 = slice_107[17:0];
assign addW_178 = concat_126 + subW_177;
assign addW_44 = slice_33 + slice_10;
assign addW_233 = add_221 + add_232;
assign subW_99 = concat_98 - concat_31;
assign slice_154 = slice_146[4:0];
assign slice_20 = slice_10[6:0];
assign concat_209 = {mul_190,slice_208};
assign lsl_75 = mulnw_74 << 10;
assign addW_130 = slice_123 + slice_108;
assign mul_51 = slice_47 * slice_50;
assign slice_240 = concat_180[31:0];
assign slice_106 = slice_105[13:7];
assign slice_161 = slice_145[8:5];
assign mul_27 = slice_20 * slice_16;
assign mulnw_216 = slice_211 * slice_198;
assign add_82 = lsl_80 + mul_81;
assign slice_137 = mul_136[9:5];
assign slice_192 = addW_186[15:0];
assign mul_113 = slice_111 * slice_112;
assign lsl_168 = add_167 << 5;
assign slice_34 = slice_14[17:0];
assign mulnw_223 = slice_193 * slice_222;
assign mulnw_89 = slice_84 * slice_54;
assign concat_144 = {addW_142,slice_143};
assign slice_10 = slice_7[31:18];
assign mul_199 = slice_197 * slice_198;
assign slice_120 = mul_113[6:0];
assign concat_175 = {addW_173,slice_174};
assign mul_230 = slice_197 * slice_226;
assign addW_96 = concat_70 + addW_95;
assign mulnw_151 = slice_129 * slice_150;
assign mul_17 = slice_12 * slice_16;
assign slice_206 = mul_199[7:0];
assign addW_127 = slice_122 + slice_105;
assign concat_182 = {concat_103,slice_181};
assign addW_48 = slice_34 + slice_15;
assign subW_237 = concat_236 - concat_103;
assign concat_103 = {addW_101,slice_102};
assign mul_158 = slice_134 * slice_154;
assign concat_24 = {mul_17,slice_23};
assign lsl_213 = mulnw_212 << 16;
assign add_79 = mulnw_76 + mulnw_78;
assign slice_134 = slice_128[4:0];
assign OUTPUT = concat_241;
    endmodule