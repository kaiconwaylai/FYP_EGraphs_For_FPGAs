//Alpha = 0.004. Cost: LUTs = 1458. DSPs = 144.  

`timescale 1ns / 1ps
    module mult(
        input[129:0] IN1,
        input[129:0] IN2,
        output[259:0] OUTPUT
    );
wire [7:0] slice_189;
wire [17:0] mul_378;
wire [27:0] add_55;
wire [16:0] slice_244;
wire [7:0] slice_110;
wire [15:0] slice_299;
wire [16:0] mul4_165;
wire [16:0] mul4_354;
wire [16:0] mul4_31;
wire [7:0] slice_220;
wire [195:0] addW_409;
wire [8:0] slice_86;
wire [64:0] slice_275;
wire [34:0] addW_141;
wire [31:0] mul_330;
wire [17:0] add_196;
wire [25:0] addW_385;
wire [16:0] mulnw_62;
wire [16:0] mul4_251;
wire [33:0] concat_117;
wire [33:0] addW_306;
wire [31:0] mul_172;
wire [8:0] slice_361;
wire [15:0] slice_38;
wire [33:0] concat_227;
wire [15:0] mul_93;
wire [8:0] slice_282;
wire [31:0] slice_148;
wire [15:0] slice_337;
wire [15:0] slice_203;
wire [16:0] mul4_392;
wire [33:0] add_69;
wire [7:0] slice_258;
wire [25:0] concat_124;
wire [32:0] slice_313;
wire [8:0] slice_179;
wire [7:0] slice_368;
wire [6:0] slice_45;
wire [7:0] slice_234;
wire [7:0] slice_100;
wire [7:0] slice_289;
wire [32:0] slice_155;
wire [8:0] slice_344;
wire [17:0] mul_21;
wire [33:0] addW_210;
wire [51:0] addW_399;
wire [63:0] mul_76;
wire [33:0] concat_265;
wire [17:0] mul_131;
wire [7:0] slice_320;
wire [27:0] add_186;
wire [33:0] concat_375;
wire [17:0] add_52;
wire [25:0] addW_241;
wire [7:0] slice_107;
wire [25:0] addW_296;
wire [7:0] slice_162;
wire [15:0] mul_351;
wire [7:0] slice_28;
wire [7:0] slice_217;
wire [132:0] concat_406;
wire [97:0] addW_272;
wire [25:0] addW_138;
wire [33:0] concat_327;
wire [16:0] mulnw_193;
wire [16:0] mul4_382;
wire [14:0] mulnw_59;
wire [7:0] slice_248;
wire [17:0] addW_114;
wire [49:0] concat_303;
wire [33:0] concat_169;
wire [7:0] slice_358;
wire [7:0] slice_35;
wire [17:0] addW_224;
wire [17:0] mul_90;
wire [65:0] addW_279;
wire [65:0] subW_145;
wire [32:0] mul4_334;
wire [32:0] slice_11;
wire [33:0] add_200;
wire [15:0] mul_389;
wire [26:0] lsl_66;
wire [33:0] concat_255;
wire [17:0] mul_121;
wire [32:0] slice_310;
wire [6:0] slice_176;
wire [7:0] slice_365;
wire [49:0] concat_42;
wire [8:0] slice_231;
wire [16:0] mul4_97;
wire [8:0] slice_286;
wire [16:0] slice_152;
wire [32:0] slice_18;
wire [63:0] mul_207;
wire [7:0] slice_396;
wire [65:0] concat_73;
wire [17:0] addW_262;
wire [25:0] addW_128;
wire [7:0] slice_317;
wire [17:0] add_183;
wire [17:0] addW_372;
wire [15:0] mulnw_49;
wire [16:0] mul4_238;
wire [16:0] slice_104;
wire [16:0] mul4_293;
wire [7:0] slice_159;
wire [17:0] mul_348;
wire [7:0] slice_25;
wire [16:0] slice_214;
wire [66:0] subW_403;
wire [68:0] concat_269;
wire [16:0] mul4_135;
wire [17:0] addW_324;
wire [14:0] mulnw_190;
wire [15:0] mul_379;
wire [33:0] add_56;
wire [50:0] concat_245;
wire [25:0] concat_111;
wire [15:0] slice_300;
wire [17:0] addW_166;
wire [16:0] mul4_355;
wire [16:0] mul4_32;
wire [25:0] concat_221;
wire [64:0] slice_410;
wire [33:0] addW_87;
wire [194:0] concat_276;
wire [51:0] addW_142;
wire [15:0] slice_331;
wire [64:0] slice_8;
wire [26:0] lsl_197;
wire [7:0] slice_386;
wire [8:0] slice_63;
wire [17:0] addW_252;
wire [16:0] slice_118;
wire [49:0] addW_307;
wire [15:0] slice_173;
wire [16:0] slice_362;
wire [31:0] mul_39;
wire [16:0] slice_228;
wire [7:0] slice_94;
wire [65:0] addW_283;
wire [129:0] concat_149;
wire [65:0] concat_338;
wire [8:0] slice_15;
wire [65:0] concat_204;
wire [16:0] mul4_393;
wire [33:0] addW_70;
wire [25:0] concat_259;
wire [16:0] mul4_125;
wire [16:0] slice_314;
wire [15:0] mulnw_180;
wire [25:0] concat_369;
wire [14:0] mulnw_46;
wire [15:0] mul_235;
wire [33:0] concat_101;
wire [15:0] mul_290;
wire [16:0] slice_156;
wire [33:0] addW_345;
wire [16:0] slice_211;
wire [16:0] slice_400;
wire [34:0] addW_266;
wire [15:0] mul_132;
wire [25:0] concat_321;
wire [33:0] add_187;
wire [16:0] slice_376;
wire [26:0] lsl_53;
wire [7:0] slice_242;
wire [7:0] slice_108;
wire [7:0] slice_297;
wire [25:0] concat_163;
wire [7:0] slice_352;
wire [25:0] concat_29;
wire [7:0] slice_218;
wire [130:0] subW_407;
wire [31:0] slice_273;
wire [7:0] slice_139;
wire [15:0] slice_328;
wire [8:0] slice_194;
wire [16:0] mul4_383;
wire [32:0] lsl_60;
wire [25:0] concat_249;
wire [25:0] addW_115;
wire [32:0] mul4_304;
wire [15:0] slice_170;
wire [33:0] concat_359;
wire [33:0] concat_36;
wire [25:0] addW_225;
wire [7:0] slice_91;
wire [32:0] slice_280;
wire [65:0] subW_146;
wire [33:0] addW_335;
wire [33:0] addW_201;
wire [7:0] slice_390;
wire [17:0] mulnw_67;
wire [17:0] mul_256;
wire [15:0] mul_122;
wire [16:0] slice_311;
wire [14:0] mulnw_177;
wire [7:0] slice_366;
wire [17:0] mul_232;
wire [17:0] addW_98;
wire [17:0] mul_287;
wire [8:0] slice_153;
wire [33:0] addW_342;
wire [16:0] slice_19;
wire [31:0] slice_208;
wire [33:0] concat_397;
wire [31:0] slice_74;
wire [25:0] addW_263;
wire [7:0] slice_129;
wire [7:0] slice_318;
wire [26:0] lsl_184;
wire [25:0] addW_373;
wire [8:0] slice_50;
wire [16:0] mul4_239;
wire [8:0] slice_105;
wire [16:0] mul4_294;
wire [7:0] slice_160;
wire [7:0] slice_349;
wire [15:0] mul_26;
wire [8:0] slice_215;
wire [99:0] addW_404;
wire [65:0] subW_270;
wire [16:0] mul4_136;
wire [25:0] addW_325;
wire [32:0] lsl_191;
wire [7:0] slice_380;
wire [6:0] slice_57;
wire [17:0] mul_246;
wire [16:0] mul4_112;
wire [31:0] mul_301;
wire [25:0] addW_167;
wire [17:0] addW_356;
wire [17:0] addW_33;
wire [16:0] mul4_222;
wire [260:0] concat_411;
wire [16:0] slice_88;
wire [16:0] slice_143;
wire [49:0] concat_332;
wire [17:0] mulnw_198;
wire [33:0] concat_387;
wire [15:0] mulnw_64;
wire [25:0] addW_253;
wire [50:0] concat_119;
wire [15:0] slice_308;
wire [49:0] concat_174;
wire [8:0] slice_363;
wire [8:0] slice_229;
wire [25:0] concat_95;
wire [32:0] slice_284;
wire [64:0] slice_150;
wire [32:0] slice_339;
wire [31:0] slice_205;
wire [17:0] addW_394;
wire [49:0] addW_71;
wire [16:0] mul4_260;
wire [16:0] mul4_126;
wire [8:0] slice_315;
wire [8:0] slice_181;
wire [16:0] mul4_370;
wire [32:0] lsl_47;
wire [7:0] slice_236;
wire [16:0] slice_102;
wire [7:0] slice_291;
wire [8:0] slice_157;
wire [16:0] slice_346;
wire [8:0] slice_212;
wire [68:0] concat_401;
wire [31:0] slice_78;
wire [51:0] addW_267;
wire [7:0] slice_133;
wire [16:0] mul4_322;
wire [6:0] slice_188;
wire [50:0] concat_377;
wire [17:0] mulnw_54;
wire [33:0] concat_243;
wire [15:0] mul_109;
wire [33:0] concat_298;
wire [16:0] mul4_164;
wire [25:0] concat_353;
wire [15:0] mul_219;
wire [130:0] subW_408;
wire [16:0] slice_85;
wire [129:0] concat_274;
wire [33:0] concat_140;
wire [15:0] slice_329;
wire [15:0] mulnw_195;
wire [17:0] addW_384;
wire [8:0] slice_61;
wire [16:0] mul4_250;
wire [7:0] slice_116;
wire [32:0] mul4_305;
wire [15:0] slice_171;
wire [16:0] slice_360;
wire [15:0] slice_37;
wire [7:0] slice_226;
wire [7:0] slice_92;
wire [16:0] slice_281;
wire [97:0] addW_147;
wire [49:0] addW_336;
wire [16:0] slice_13;
wire [49:0] addW_202;
wire [25:0] concat_391;
wire [27:0] add_68;
wire [15:0] mul_257;
wire [7:0] slice_123;
wire [8:0] slice_312;
wire [32:0] lsl_178;
wire [15:0] mul_367;
wire [7:0] slice_44;
wire [7:0] slice_233;
wire [25:0] addW_99;
wire [7:0] slice_288;
wire [64:0] slice_154;
wire [16:0] slice_343;
wire [8:0] slice_20;
wire [97:0] concat_209;
wire [34:0] addW_398;
wire [31:0] slice_75;
wire [7:0] slice_264;
wire [33:0] concat_130;
wire [15:0] mul_319;
wire [17:0] mulnw_185;
wire [7:0] slice_374;
wire [16:0] mulnw_51;
wire [17:0] addW_240;
wire [17:0] mul_106;
wire [17:0] addW_295;
wire [15:0] mul_161;
wire [7:0] slice_350;
wire [17:0] mul_216;
wire [32:0] slice_405;
wire [33:0] addW_82;
wire [65:0] subW_271;
wire [17:0] addW_137;
wire [7:0] slice_326;
wire [8:0] slice_192;
wire [25:0] concat_381;
wire [7:0] slice_58;
wire [15:0] mul_247;
wire [16:0] mul4_113;
wire [15:0] slice_302;
wire [7:0] slice_168;
wire [25:0] addW_357;
wire [25:0] addW_34;
wire [16:0] mul4_223;
wire [8:0] slice_89;
wire [68:0] concat_144;
wire [32:0] mul4_333;
wire [27:0] add_199;
wire [17:0] mul_388;
wire [17:0] add_65;
wire [7:0] slice_254;
wire [65:0] concat_309;
wire [7:0] slice_175;
wire [17:0] mul_364;
wire [15:0] slice_41;
wire [16:0] slice_230;
wire [16:0] mul4_96;
wire [16:0] slice_285;
wire [32:0] slice_151;
wire [98:0] concat_340;
wire [64:0] slice_17;
wire [31:0] slice_206;
wire [25:0] addW_395;
wire [15:0] slice_72;
wire [16:0] mul4_261;
wire [17:0] addW_127;
wire [17:0] mul_316;
wire [16:0] mulnw_182;
wire [16:0] mul4_371;
wire [8:0] slice_48;
wire [25:0] concat_237;
wire [8:0] slice_103;
wire [25:0] concat_292;
wire [17:0] mul_158;
wire [8:0] slice_347;
wire [7:0] slice_24;
wire [33:0] addW_213;
wire [66:0] subW_402;
wire [97:0] concat_79;
wire [16:0] slice_268;
wire [25:0] concat_134;
wire [16:0] mul4_323;
assign slice_189 = slice_156[16:9];
assign mul_378 = slice_344 * slice_363;
assign add_55 = lsl_53 + mulnw_54;
assign slice_244 = concat_243[33:17];
assign slice_110 = mul_109[15:8];
assign slice_299 = slice_280[15:0];
assign mul4_165 = slice_159 * slice_157;
assign mul4_354 = slice_344 * slice_350;
assign mul4_31 = slice_15 * slice_25;
assign slice_220 = mul_219[15:8];
assign addW_409 = concat_276 + subW_408;
assign slice_86 = slice_85[16:8];
assign slice_275 = concat_274[129:65];
assign addW_141 = concat_130 + concat_140;
assign mul_330 = slice_328 * slice_329;
assign add_196 = mulnw_193 + mulnw_195;
assign addW_385 = concat_381 + addW_384;
assign mulnw_62 = slice_61 * slice_58;
assign mul4_251 = slice_217 * slice_231;
assign concat_117 = {addW_115,slice_116};
assign addW_306 = mul4_304 + mul4_305;
assign mul_172 = slice_170 * slice_171;
assign slice_361 = slice_360[16:8];
assign slice_38 = slice_18[15:0];
assign concat_227 = {addW_225,slice_226};
assign mul_93 = slice_91 * slice_92;
assign slice_282 = slice_281[16:8];
assign slice_148 = mul_76[31:0];
assign slice_337 = mul_330[15:0];
assign slice_203 = mul_172[15:0];
assign mul4_392 = slice_361 * slice_350;
assign add_69 = lsl_60 + add_68;
assign slice_258 = mul_257[15:8];
assign concat_124 = {mul_121,slice_123};
assign slice_313 = addW_283[32:0];
assign slice_179 = slice_152[8:0];
assign slice_368 = mul_367[15:8];
assign slice_45 = slice_38[15:9];
assign slice_234 = slice_230[7:0];
assign slice_100 = mul_93[7:0];
assign slice_289 = slice_285[7:0];
assign slice_155 = slice_154[64:32];
assign slice_344 = slice_343[16:8];
assign mul_21 = slice_15 * slice_20;
assign addW_210 = slice_205 + slice_151;
assign addW_399 = concat_377 + addW_398;
assign mul_76 = slice_74 * slice_75;
assign concat_265 = {addW_263,slice_264};
assign mul_131 = slice_103 * slice_89;
assign slice_320 = mul_319[15:8];
assign add_186 = lsl_184 + mulnw_185;
assign concat_375 = {addW_373,slice_374};
assign add_52 = mulnw_49 + mulnw_51;
assign addW_241 = concat_237 + addW_240;
assign slice_107 = slice_102[7:0];
assign addW_296 = concat_292 + addW_295;
assign slice_162 = mul_161[15:8];
assign mul_351 = slice_349 * slice_350;
assign slice_28 = mul_26[15:8];
assign slice_217 = slice_211[7:0];
assign concat_406 = {addW_404,slice_405};
assign addW_272 = concat_209 + subW_271;
assign addW_138 = concat_134 + addW_137;
assign concat_327 = {addW_325,slice_326};
assign mulnw_193 = slice_192 * slice_189;
assign mul4_382 = slice_344 * slice_366;
assign mulnw_59 = slice_57 * slice_58;
assign slice_248 = mul_247[15:8];
assign addW_114 = mul4_112 + mul4_113;
assign concat_303 = {concat_298,slice_302};
assign concat_169 = {addW_167,slice_168};
assign slice_358 = mul_351[7:0];
assign slice_35 = mul_26[7:0];
assign addW_224 = mul4_222 + mul4_223;
assign mul_90 = slice_86 * slice_89;
assign addW_279 = slice_150 + slice_8;
assign subW_145 = concat_144 - concat_73;
assign mul4_334 = slice_328 * slice_314;
assign slice_11 = slice_8[64:32];
assign add_200 = lsl_191 + add_199;
assign mul_389 = slice_365 * slice_350;
assign lsl_66 = add_65 << 9;
assign concat_255 = {addW_253,slice_254};
assign mul_121 = slice_86 * slice_105;
assign slice_310 = addW_279[32:0];
assign slice_176 = slice_171[15:9];
assign slice_365 = slice_360[7:0];
assign concat_42 = {concat_36,slice_41};
assign slice_231 = slice_230[16:8];
assign mul4_97 = slice_91 * slice_89;
assign slice_286 = slice_285[16:8];
assign slice_152 = slice_151[32:16];
assign slice_18 = slice_17[64:32];
assign mul_207 = slice_205 * slice_206;
assign slice_396 = mul_389[7:0];
assign concat_73 = {addW_71,slice_72};
assign addW_262 = mul4_260 + mul4_261;
assign addW_128 = concat_124 + addW_127;
assign slice_317 = slice_311[7:0];
assign add_183 = mulnw_180 + mulnw_182;
assign addW_372 = mul4_370 + mul4_371;
assign mulnw_49 = slice_48 * slice_45;
assign mul4_238 = slice_229 * slice_234;
assign slice_104 = addW_87[16:0];
assign mul4_293 = slice_282 * slice_289;
assign slice_159 = slice_152[7:0];
assign mul_348 = slice_344 * slice_347;
assign slice_25 = slice_19[7:0];
assign slice_214 = addW_213[33:17];
assign subW_403 = subW_402 - concat_338;
assign concat_269 = {addW_267,slice_268};
assign mul4_135 = slice_103 * slice_92;
assign addW_324 = mul4_322 + mul4_323;
assign mulnw_190 = slice_188 * slice_189;
assign mul_379 = slice_349 * slice_366;
assign add_56 = lsl_47 + add_55;
assign concat_245 = {concat_227,slice_244};
assign concat_111 = {mul_106,slice_110};
assign slice_300 = slice_284[15:0];
assign addW_166 = mul4_164 + mul4_165;
assign mul4_355 = slice_349 * slice_347;
assign mul4_32 = slice_24 * slice_20;
assign concat_221 = {mul_216,slice_220};
assign slice_410 = concat_274[64:0];
assign addW_87 = slice_75 + slice_18;
assign concat_276 = {concat_149,slice_275};
assign addW_142 = concat_119 + addW_141;
assign slice_331 = mul_330[31:16];
assign slice_8 = IN1[129:65];
assign lsl_197 = add_196 << 9;
assign slice_386 = mul_379[7:0];
assign slice_63 = slice_19[8:0];
assign addW_252 = mul4_250 + mul4_251;
assign slice_118 = concat_117[33:17];
assign addW_307 = concat_303 + addW_306;
assign slice_173 = mul_172[31:16];
assign slice_362 = addW_345[16:0];
assign mul_39 = slice_37 * slice_38;
assign slice_228 = addW_210[16:0];
assign slice_94 = mul_93[15:8];
assign addW_283 = slice_154 + slice_17;
assign concat_149 = {addW_147,slice_148};
assign concat_338 = {addW_336,slice_337};
assign slice_15 = slice_13[16:8];
assign concat_204 = {addW_202,slice_203};
assign mul4_393 = slice_365 * slice_347;
assign addW_70 = add_56 + add_69;
assign concat_259 = {mul_256,slice_258};
assign mul4_125 = slice_86 * slice_108;
assign slice_314 = slice_313[32:16];
assign mulnw_180 = slice_179 * slice_176;
assign concat_369 = {mul_364,slice_368};
assign mulnw_46 = slice_44 * slice_45;
assign mul_235 = slice_233 * slice_234;
assign concat_101 = {addW_99,slice_100};
assign mul_290 = slice_288 * slice_289;
assign slice_156 = slice_155[32:16];
assign addW_345 = slice_313 + slice_284;
assign slice_211 = addW_210[33:17];
assign slice_400 = concat_375[16:0];
assign addW_266 = concat_255 + concat_265;
assign mul_132 = slice_107 * slice_92;
assign concat_321 = {mul_316,slice_320};
assign add_187 = lsl_178 + add_186;
assign slice_376 = concat_375[33:17];
assign lsl_53 = add_52 << 9;
assign slice_242 = mul_235[7:0];
assign slice_108 = slice_104[7:0];
assign slice_297 = mul_290[7:0];
assign concat_163 = {mul_158,slice_162};
assign slice_352 = mul_351[15:8];
assign concat_29 = {mul_21,slice_28};
assign slice_218 = slice_214[7:0];
assign subW_407 = concat_406 - concat_149;
assign slice_273 = mul_207[31:0];
assign slice_139 = mul_132[7:0];
assign slice_328 = slice_310[15:0];
assign slice_194 = slice_156[8:0];
assign mul4_383 = slice_349 * slice_363;
assign lsl_60 = mulnw_59 << 18;
assign concat_249 = {mul_246,slice_248};
assign addW_115 = concat_111 + addW_114;
assign mul4_304 = slice_281 * slice_300;
assign slice_170 = slice_151[15:0];
assign concat_359 = {addW_357,slice_358};
assign concat_36 = {addW_34,slice_35};
assign addW_225 = concat_221 + addW_224;
assign slice_91 = slice_85[7:0];
assign slice_280 = addW_279[65:33];
assign subW_146 = subW_145 - mul_76;
assign addW_335 = mul4_333 + mul4_334;
assign addW_201 = add_187 + add_200;
assign slice_390 = mul_389[15:8];
assign mulnw_67 = slice_61 * slice_63;
assign mul_256 = slice_229 * slice_215;
assign mul_122 = slice_91 * slice_108;
assign slice_311 = slice_310[32:16];
assign mulnw_177 = slice_175 * slice_176;
assign slice_366 = slice_362[7:0];
assign mul_232 = slice_229 * slice_231;
assign addW_98 = mul4_96 + mul4_97;
assign mul_287 = slice_282 * slice_286;
assign slice_153 = slice_152[16:8];
assign addW_342 = slice_310 + slice_280;
assign slice_19 = slice_18[32:16];
assign slice_208 = mul_207[63:32];
assign concat_397 = {addW_395,slice_396};
assign slice_74 = slice_8[31:0];
assign addW_263 = concat_259 + addW_262;
assign slice_129 = mul_122[7:0];
assign slice_318 = slice_314[7:0];
assign lsl_184 = add_183 << 9;
assign addW_373 = concat_369 + addW_372;
assign slice_50 = slice_38[8:0];
assign mul4_239 = slice_233 * slice_231;
assign slice_105 = slice_104[16:8];
assign mul4_294 = slice_288 * slice_286;
assign slice_160 = slice_156[7:0];
assign slice_349 = slice_343[7:0];
assign mul_26 = slice_24 * slice_25;
assign slice_215 = slice_214[16:8];
assign addW_404 = concat_340 + subW_403;
assign subW_270 = concat_269 - concat_204;
assign mul4_136 = slice_107 * slice_89;
assign addW_325 = concat_321 + addW_324;
assign lsl_191 = mulnw_190 << 18;
assign slice_380 = mul_379[15:8];
assign slice_57 = slice_37[15:9];
assign mul_246 = slice_212 * slice_231;
assign mul4_112 = slice_103 * slice_108;
assign mul_301 = slice_299 * slice_300;
assign addW_167 = concat_163 + addW_166;
assign addW_356 = mul4_354 + mul4_355;
assign addW_33 = mul4_31 + mul4_32;
assign mul4_222 = slice_212 * slice_218;
assign concat_411 = {addW_409,slice_410};
assign slice_88 = addW_87[33:17];
assign slice_143 = concat_117[16:0];
assign concat_332 = {concat_327,slice_331};
assign mulnw_198 = slice_192 * slice_194;
assign concat_387 = {addW_385,slice_386};
assign mulnw_64 = slice_57 * slice_63;
assign addW_253 = concat_249 + addW_252;
assign concat_119 = {concat_101,slice_118};
assign slice_308 = mul_301[15:0];
assign concat_174 = {concat_169,slice_173};
assign slice_363 = slice_362[16:8];
assign slice_229 = slice_228[16:8];
assign concat_95 = {mul_90,slice_94};
assign slice_284 = addW_283[65:33];
assign slice_150 = IN1[64:0];
assign slice_339 = concat_338[65:33];
assign slice_205 = slice_150[31:0];
assign addW_394 = mul4_392 + mul4_393;
assign addW_71 = concat_42 + addW_70;
assign mul4_260 = slice_229 * slice_218;
assign mul4_126 = slice_91 * slice_105;
assign slice_315 = slice_314[16:8];
assign slice_181 = slice_171[8:0];
assign mul4_370 = slice_361 * slice_366;
assign lsl_47 = mulnw_46 << 18;
assign slice_236 = mul_235[15:8];
assign slice_102 = addW_82[16:0];
assign slice_291 = mul_290[15:8];
assign slice_157 = slice_156[16:8];
assign slice_346 = addW_345[33:17];
assign slice_212 = slice_211[16:8];
assign concat_401 = {addW_399,slice_400};
assign slice_78 = mul_76[63:32];
assign addW_267 = concat_245 + addW_266;
assign slice_133 = mul_132[15:8];
assign mul4_322 = slice_312 * slice_318;
assign slice_188 = slice_170[15:9];
assign concat_377 = {concat_359,slice_376};
assign mulnw_54 = slice_48 * slice_50;
assign concat_243 = {addW_241,slice_242};
assign mul_109 = slice_107 * slice_108;
assign concat_298 = {addW_296,slice_297};
assign mul4_164 = slice_153 * slice_160;
assign concat_353 = {mul_348,slice_352};
assign mul_219 = slice_217 * slice_218;
assign subW_408 = subW_407 - concat_274;
assign slice_85 = addW_82[33:17];
assign concat_274 = {addW_272,slice_273};
assign concat_140 = {addW_138,slice_139};
assign slice_329 = slice_313[15:0];
assign mulnw_195 = slice_188 * slice_194;
assign addW_384 = mul4_382 + mul4_383;
assign slice_61 = slice_37[8:0];
assign mul4_250 = slice_212 * slice_234;
assign slice_116 = mul_109[7:0];
assign mul4_305 = slice_299 * slice_285;
assign slice_171 = slice_155[15:0];
assign slice_360 = addW_342[16:0];
assign slice_37 = slice_11[15:0];
assign slice_226 = mul_219[7:0];
assign slice_92 = slice_88[7:0];
assign slice_281 = slice_280[32:16];
assign addW_147 = concat_79 + subW_146;
assign addW_336 = concat_332 + addW_335;
assign slice_13 = slice_11[32:16];
assign addW_202 = concat_174 + addW_201;
assign concat_391 = {mul_388,slice_390};
assign add_68 = lsl_66 + mulnw_67;
assign mul_257 = slice_233 * slice_218;
assign slice_123 = mul_122[15:8];
assign slice_312 = slice_311[16:8];
assign lsl_178 = mulnw_177 << 18;
assign mul_367 = slice_365 * slice_366;
assign slice_44 = slice_13[16:9];
assign slice_233 = slice_228[7:0];
assign addW_99 = concat_95 + addW_98;
assign slice_288 = slice_281[7:0];
assign slice_154 = IN2[64:0];
assign slice_343 = addW_342[33:17];
assign slice_20 = slice_19[16:8];
assign concat_209 = {concat_204,slice_208};
assign addW_398 = concat_387 + concat_397;
assign slice_75 = slice_17[31:0];
assign slice_264 = mul_257[7:0];
assign concat_130 = {addW_128,slice_129};
assign mul_319 = slice_317 * slice_318;
assign mulnw_185 = slice_179 * slice_181;
assign slice_374 = mul_367[7:0];
assign mulnw_51 = slice_44 * slice_50;
assign addW_240 = mul4_238 + mul4_239;
assign mul_106 = slice_103 * slice_105;
assign addW_295 = mul4_293 + mul4_294;
assign mul_161 = slice_159 * slice_160;
assign slice_350 = slice_346[7:0];
assign mul_216 = slice_212 * slice_215;
assign slice_405 = concat_338[32:0];
assign addW_82 = slice_74 + slice_11;
assign subW_271 = subW_270 - mul_207;
assign addW_137 = mul4_135 + mul4_136;
assign slice_326 = mul_319[7:0];
assign slice_192 = slice_170[8:0];
assign concat_381 = {mul_378,slice_380};
assign slice_58 = slice_19[16:9];
assign mul_247 = slice_217 * slice_234;
assign mul4_113 = slice_107 * slice_105;
assign slice_302 = mul_301[31:16];
assign slice_168 = mul_161[7:0];
assign addW_357 = concat_353 + addW_356;
assign addW_34 = concat_29 + addW_33;
assign mul4_223 = slice_217 * slice_215;
assign slice_89 = slice_88[16:8];
assign concat_144 = {addW_142,slice_143};
assign mul4_333 = slice_311 * slice_329;
assign add_199 = lsl_197 + mulnw_198;
assign mul_388 = slice_361 * slice_347;
assign add_65 = mulnw_62 + mulnw_64;
assign slice_254 = mul_247[7:0];
assign concat_309 = {addW_307,slice_308};
assign slice_175 = slice_152[16:9];
assign mul_364 = slice_361 * slice_363;
assign slice_41 = mul_39[31:16];
assign slice_230 = addW_213[16:0];
assign mul4_96 = slice_86 * slice_92;
assign slice_285 = slice_284[32:16];
assign slice_151 = slice_150[64:32];
assign concat_340 = {concat_309,slice_339};
assign slice_17 = IN2[129:65];
assign slice_206 = slice_154[31:0];
assign addW_395 = concat_391 + addW_394;
assign slice_72 = mul_39[15:0];
assign mul4_261 = slice_233 * slice_215;
assign addW_127 = mul4_125 + mul4_126;
assign mul_316 = slice_312 * slice_315;
assign mulnw_182 = slice_175 * slice_181;
assign mul4_371 = slice_365 * slice_363;
assign slice_48 = slice_13[8:0];
assign concat_237 = {mul_232,slice_236};
assign slice_103 = slice_102[16:8];
assign concat_292 = {mul_287,slice_291};
assign mul_158 = slice_153 * slice_157;
assign slice_347 = slice_346[16:8];
assign slice_24 = slice_13[7:0];
assign addW_213 = slice_206 + slice_155;
assign subW_402 = concat_401 - concat_309;
assign concat_79 = {concat_73,slice_78};
assign slice_268 = concat_243[16:0];
assign concat_134 = {mul_131,slice_133};
assign mul4_323 = slice_317 * slice_315;
assign OUTPUT = concat_411;
    endmodule