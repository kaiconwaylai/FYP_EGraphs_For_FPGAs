//Alpha = 0.005. Cost: LUTs = 3483. DSPs = 0.  

`timescale 1ns / 1ps
    module mult(
        input[255:0] IN1,
        input[255:0] IN2,
        output[511:0] OUTPUT
    );
wire [26:0] add_189;
wire [67:0] subW_378;
wire [16:0] slice_567;
wire [7:0] slice_756;
wire [67:0] subW_110;
wire [13:0] slice_299;
wire [7:0] slice_488;
wire [17:0] slice_677;
wire [45:0] concat_31;
wire [7:0] slice_220;
wire [17:0] slice_409;
wire [15:0] mulnw_598;
wire [15:0] slice_787;
wire [17:0] slice_141;
wire [39:0] mul_330;
wire [35:0] mul_519;
wire [16:0] mulnw_708;
wire [17:0] slice_251;
wire [16:0] mulnw_440;
wire [15:0] slice_629;
wire [34:0] addW_818;
wire [16:0] mulnw_172;
wire [7:0] slice_361;
wire [70:0] subW_550;
wire [7:0] slice_93;
wire [41:0] subW_282;
wire [32:0] slice_471;
wire [35:0] mul_660;
wire [135:0] subW_849;
wire [31:0] slice_14;
wire [35:0] mul_392;
wire [32:0] lsl_581;
wire [16:0] mulnw_770;
wire [35:0] mul_124;
wire [40:0] subW_313;
wire [15:0] mulnw_502;
wire [33:0] addW_691;
wire [13:0] slice_45;
wire [16:0] mulnw_234;
wire [33:0] addW_423;
wire [27:0] mul_612;
wire [25:0] lsl_801;
wire [33:0] addW_155;
wire [15:0] slice_344;
wire [15:0] slice_533;
wire [17:0] add_722;
wire [49:0] concat_76;
wire [98:0] concat_265;
wire [17:0] add_454;
wire [51:0] addW_643;
wire [35:0] mul_832;
wire [17:0] add_186;
wire [50:0] addW_375;
wire [129:0] addW_564;
wire [7:0] slice_753;
wire [50:0] addW_107;
wire [127:0] slice_296;
wire [32:0] lsl_485;
wire [13:0] slice_674;
wire [35:0] mul_28;
wire [7:0] slice_217;
wire [13:0] slice_406;
wire [7:0] slice_595;
wire [32:0] slice_784;
wire [13:0] slice_138;
wire [45:0] concat_327;
wire [27:0] mul_516;
wire [7:0] slice_705;
wire [65:0] concat_59;
wire [31:0] slice_248;
wire [7:0] slice_437;
wire [31:0] slice_626;
wire [15:0] mul_815;
wire [7:0] slice_169;
wire [15:0] mul_358;
wire [51:0] addW_547;
wire [63:0] slice_736;
wire [15:0] mul_90;
wire [19:0] addW_279;
wire [63:0] slice_468;
wire [27:0] mul_657;
wire [32:0] slice_846;
wire [63:0] slice_11;
wire [63:0] slice_200;
wire [27:0] mul_389;
wire [8:0] slice_578;
wire [16:0] mulnw_767;
wire [27:0] mul_121;
wire [19:0] addW_310;
wire [7:0] slice_499;
wire [65:0] concat_688;
wire [31:0] slice_42;
wire [16:0] mulnw_231;
wire [65:0] concat_420;
wire [13:0] slice_609;
wire [7:0] slice_798;
wire [65:0] concat_152;
wire [16:0] slice_341;
wire [31:0] slice_530;
wire [16:0] mulnw_719;
wire [15:0] slice_73;
wire [17:0] slice_262;
wire [16:0] mulnw_451;
wire [39:0] mul_640;
wire [31:0] mul_829;
wire [16:0] mulnw_183;
wire [26:0] add_372;
wire [387:0] concat_561;
wire [15:0] slice_750;
wire [26:0] add_104;
wire [195:0] addW_293;
wire [8:0] slice_482;
wire [31:0] slice_671;
wire [15:0] slice_214;
wire [31:0] slice_403;
wire [8:0] slice_592;
wire [66:0] concat_781;
wire [31:0] slice_135;
wire [17:0] slice_324;
wire [13:0] slice_513;
wire [7:0] slice_702;
wire [41:0] subW_56;
wire [66:0] concat_245;
wire [7:0] slice_434;
wire [47:0] addW_623;
wire [15:0] mulnw_812;
wire [7:0] slice_166;
wire [16:0] mulnw_355;
wire [39:0] mul_544;
wire [98:0] addW_733;
wire [16:0] mulnw_87;
wire [17:0] slice_276;
wire [98:0] addW_465;
wire [63:0] slice_654;
wire [70:0] subW_843;
wire [127:0] slice_8;
wire [98:0] addW_197;
wire [63:0] slice_386;
wire [31:0] mul_575;
wire [33:0] add_764;
wire [63:0] slice_118;
wire [35:0] mul_307;
wire [8:0] slice_496;
wire [41:0] subW_685;
wire [47:0] addW_39;
wire [33:0] add_228;
wire [41:0] subW_417;
wire [15:0] slice_606;
wire [32:0] lsl_795;
wire [41:0] subW_149;
wire [33:0] addW_338;
wire [47:0] addW_527;
wire [16:0] mulnw_716;
wire [33:0] mul_70;
wire [40:0] subW_259;
wire [16:0] mulnw_448;
wire [49:0] concat_637;
wire [15:0] slice_826;
wire [16:0] mulnw_180;
wire [17:0] add_369;
wire [63:0] slice_558;
wire [15:0] slice_747;
wire [17:0] add_101;
wire [131:0] concat_290;
wire [31:0] mul_479;
wire [47:0] addW_668;
wire [516:0] concat_857;
wire [13:0] slice_22;
wire [15:0] slice_211;
wire [47:0] addW_400;
wire [26:0] add_589;
wire [34:0] addW_778;
wire [47:0] addW_132;
wire [13:0] slice_321;
wire [15:0] slice_510;
wire [15:0] slice_699;
wire [19:0] addW_53;
wire [34:0] addW_242;
wire [15:0] slice_431;
wire [39:0] mul_620;
wire [7:0] slice_809;
wire [15:0] slice_163;
wire [7:0] slice_352;
wire [49:0] concat_541;
wire [66:0] concat_730;
wire [7:0] slice_84;
wire [17:0] slice_273;
wire [66:0] concat_462;
wire [63:0] slice_651;
wire [51:0] addW_840;
wire [66:0] concat_194;
wire [63:0] slice_383;
wire [33:0] mul_572;
wire [25:0] lsl_761;
wire [63:0] slice_115;
wire [27:0] mul_304;
wire [26:0] add_493;
wire [19:0] addW_682;
wire [39:0] mul_36;
wire [25:0] lsl_225;
wire [19:0] addW_414;
wire [33:0] add_603;
wire [8:0] slice_792;
wire [19:0] addW_146;
wire [65:0] concat_335;
wire [39:0] mul_524;
wire [33:0] add_713;
wire [16:0] slice_67;
wire [19:0] addW_256;
wire [33:0] add_445;
wire [17:0] slice_634;
wire [99:0] concat_823;
wire [33:0] add_177;
wire [16:0] mulnw_366;
wire [132:0] subW_555;
wire [32:0] slice_744;
wire [16:0] mulnw_98;
wire [71:0] subW_287;
wire [33:0] mul_476;
wire [39:0] mul_665;
wire [262:0] subW_854;
wire [127:0] slice_19;
wire [32:0] slice_208;
wire [39:0] mul_397;
wire [17:0] add_586;
wire [15:0] mul_775;
wire [39:0] mul_129;
wire [31:0] slice_318;
wire [33:0] add_507;
wire [15:0] slice_696;
wire [17:0] slice_50;
wire [15:0] mul_239;
wire [15:0] slice_428;
wire [45:0] concat_617;
wire [8:0] slice_806;
wire [15:0] slice_160;
wire [7:0] slice_349;
wire [17:0] slice_538;
wire [34:0] addW_727;
wire [16:0] mulnw_81;
wire [34:0] addW_270;
wire [34:0] addW_459;
wire [99:0] addW_648;
wire [39:0] mul_837;
wire [34:0] addW_191;
wire [98:0] addW_380;
wire [64:0] slice_569;
wire [7:0] slice_758;
wire [98:0] addW_112;
wire [63:0] slice_301;
wire [17:0] add_490;
wire [17:0] slice_679;
wire [7:0] slice_222;
wire [17:0] slice_411;
wire [25:0] lsl_600;
wire [31:0] mul_789;
wire [17:0] slice_143;
wire [41:0] subW_332;
wire [45:0] concat_521;
wire [25:0] lsl_710;
wire [35:0] mul_253;
wire [25:0] lsl_442;
wire [15:0] slice_631;
wire [15:0] slice_820;
wire [25:0] lsl_174;
wire [16:0] mulnw_363;
wire [99:0] addW_552;
wire [32:0] slice_741;
wire [16:0] mulnw_95;
wire [17:0] slice_284;
wire [65:0] addW_473;
wire [45:0] concat_662;
wire [63:0] slice_851;
wire [32:0] slice_205;
wire [45:0] concat_394;
wire [15:0] mulnw_583;
wire [15:0] mulnw_772;
wire [45:0] concat_126;
wire [47:0] addW_315;
wire [25:0] lsl_504;
wire [33:0] addW_693;
wire [17:0] slice_47;
wire [15:0] mulnw_236;
wire [33:0] addW_425;
wire [17:0] slice_614;
wire [26:0] add_803;
wire [33:0] addW_157;
wire [15:0] slice_346;
wire [15:0] slice_535;
wire [15:0] mul_724;
wire [15:0] mul_456;
wire [69:0] concat_645;
wire [49:0] concat_834;
wire [15:0] mul_188;
wire [66:0] concat_377;
wire [32:0] slice_566;
wire [32:0] lsl_755;
wire [66:0] concat_109;
wire [31:0] slice_298;
wire [15:0] mulnw_487;
wire [17:0] slice_676;
wire [17:0] slice_30;
wire [32:0] lsl_219;
wire [17:0] slice_408;
wire [7:0] slice_597;
wire [33:0] mul_786;
wire [17:0] slice_140;
wire [19:0] addW_329;
wire [17:0] slice_518;
wire [7:0] slice_707;
wire [97:0] concat_61;
wire [27:0] mul_250;
wire [7:0] slice_439;
wire [34:0] addW_628;
wire [33:0] add_817;
wire [7:0] slice_171;
wire [33:0] add_360;
wire [69:0] concat_549;
wire [33:0] add_92;
wire [40:0] subW_281;
wire [65:0] addW_470;
wire [17:0] slice_659;
wire [134:0] subW_848;
wire [17:0] slice_391;
wire [16:0] mulnw_580;
wire [7:0] slice_769;
wire [17:0] slice_123;
wire [39:0] mul_312;
wire [7:0] slice_501;
wire [97:0] concat_690;
wire [31:0] slice_44;
wire [7:0] slice_233;
wire [97:0] concat_422;
wire [13:0] slice_611;
wire [17:0] add_800;
wire [97:0] concat_154;
wire [15:0] slice_343;
wire [34:0] addW_532;
wire [15:0] mulnw_721;
wire [15:0] slice_75;
wire [31:0] slice_264;
wire [15:0] mulnw_453;
wire [41:0] subW_642;
wire [17:0] slice_831;
wire [15:0] mulnw_185;
wire [34:0] addW_374;
wire [8:0] slice_752;
wire [34:0] addW_106;
wire [259:0] concat_295;
wire [16:0] mulnw_484;
wire [31:0] slice_673;
wire [17:0] slice_27;
wire [8:0] slice_216;
wire [31:0] slice_405;
wire [32:0] lsl_594;
wire [16:0] slice_783;
wire [31:0] slice_137;
wire [17:0] slice_326;
wire [13:0] slice_515;
wire [32:0] lsl_704;
wire [17:0] slice_58;
wire [13:0] slice_247;
wire [32:0] lsl_436;
wire [65:0] concat_625;
wire [25:0] lsl_814;
wire [32:0] lsl_168;
wire [25:0] lsl_357;
wire [41:0] subW_546;
wire [130:0] concat_735;
wire [25:0] lsl_89;
wire [19:0] addW_278;
wire [130:0] concat_467;
wire [13:0] slice_656;
wire [100:0] addW_845;
wire [130:0] concat_199;
wire [13:0] slice_388;
wire [49:0] concat_577;
wire [8:0] slice_766;
wire [13:0] slice_120;
wire [45:0] concat_309;
wire [32:0] lsl_498;
wire [17:0] slice_687;
wire [65:0] concat_41;
wire [8:0] slice_230;
wire [17:0] slice_419;
wire [31:0] slice_608;
wire [15:0] mulnw_797;
wire [17:0] slice_151;
wire [33:0] addW_340;
wire [65:0] concat_529;
wire [7:0] slice_718;
wire [15:0] slice_72;
wire [47:0] addW_261;
wire [7:0] slice_450;
wire [19:0] addW_639;
wire [15:0] slice_828;
wire [7:0] slice_182;
wire [15:0] mul_371;
wire [127:0] slice_560;
wire [31:0] mul_749;
wire [15:0] mul_103;
wire [133:0] subW_292;
wire [49:0] concat_481;
wire [65:0] concat_670;
wire [31:0] mul_213;
wire [65:0] concat_402;
wire [7:0] slice_591;
wire [15:0] slice_780;
wire [65:0] concat_134;
wire [17:0] slice_323;
wire [31:0] slice_512;
wire [8:0] slice_701;
wire [40:0] subW_55;
wire [15:0] slice_244;
wire [8:0] slice_433;
wire [41:0] subW_622;
wire [7:0] slice_811;
wire [8:0] slice_165;
wire [7:0] slice_354;
wire [19:0] addW_543;
wire [68:0] subW_732;
wire [7:0] slice_86;
wire [35:0] mul_275;
wire [68:0] subW_464;
wire [13:0] slice_653;
wire [69:0] concat_842;
wire [68:0] subW_196;
wire [13:0] slice_385;
wire [15:0] slice_574;
wire [26:0] add_763;
wire [13:0] slice_117;
wire [17:0] slice_306;
wire [7:0] slice_495;
wire [40:0] subW_684;
wire [41:0] subW_38;
wire [26:0] add_227;
wire [40:0] subW_416;
wire [50:0] addW_605;
wire [16:0] mulnw_794;
wire [40:0] subW_148;
wire [97:0] concat_337;
wire [41:0] subW_526;
wire [8:0] slice_715;
wire [16:0] slice_69;
wire [39:0] mul_258;
wire [8:0] slice_447;
wire [17:0] slice_636;
wire [34:0] addW_825;
wire [8:0] slice_179;
wire [15:0] mulnw_368;
wire [195:0] addW_557;
wire [33:0] mul_746;
wire [15:0] mulnw_100;
wire [31:0] slice_289;
wire [15:0] slice_478;
wire [41:0] subW_667;
wire [127:0] slice_856;
wire [31:0] slice_21;
wire [33:0] mul_210;
wire [41:0] subW_399;
wire [15:0] mul_588;
wire [33:0] add_777;
wire [41:0] subW_131;
wire [31:0] slice_320;
wire [50:0] addW_509;
wire [31:0] mul_698;
wire [19:0] addW_52;
wire [33:0] add_241;
wire [31:0] mul_430;
wire [19:0] addW_619;
wire [32:0] lsl_808;
wire [31:0] mul_162;
wire [32:0] lsl_351;
wire [17:0] slice_540;
wire [15:0] slice_729;
wire [31:0] mul_272;
wire [15:0] slice_461;
wire [131:0] concat_650;
wire [41:0] subW_839;
wire [15:0] slice_193;
wire [130:0] concat_382;
wire [16:0] slice_571;
wire [17:0] add_760;
wire [130:0] concat_114;
wire [13:0] slice_303;
wire [15:0] mul_492;
wire [19:0] addW_681;
wire [19:0] addW_35;
wire [17:0] add_224;
wire [19:0] addW_413;
wire [26:0] add_602;
wire [49:0] concat_791;
wire [19:0] addW_145;
wire [17:0] slice_334;
wire [19:0] addW_523;
wire [26:0] add_712;
wire [45:0] concat_255;
wire [26:0] add_444;
wire [17:0] slice_633;
wire [32:0] slice_822;
wire [26:0] add_176;
wire [7:0] slice_365;
wire [131:0] concat_554;
wire [66:0] addW_743;
wire [7:0] slice_97;
wire [70:0] subW_286;
wire [16:0] slice_475;
wire [19:0] addW_664;
wire [261:0] subW_853;
wire [65:0] addW_207;
wire [19:0] addW_396;
wire [16:0] mulnw_585;
wire [25:0] lsl_774;
wire [19:0] addW_128;
wire [65:0] concat_317;
wire [26:0] add_506;
wire [33:0] mul_695;
wire [35:0] mul_49;
wire [25:0] lsl_238;
wire [33:0] mul_427;
wire [17:0] slice_616;
wire [7:0] slice_805;
wire [33:0] mul_159;
wire [8:0] slice_348;
wire [17:0] slice_537;
wire [33:0] add_726;
wire [7:0] slice_80;
wire [15:0] slice_269;
wire [33:0] add_458;
wire [71:0] subW_647;
wire [19:0] addW_836;
wire [33:0] add_190;
wire [68:0] subW_379;
wire [129:0] addW_568;
wire [15:0] mulnw_757;
wire [68:0] subW_111;
wire [127:0] slice_300;
wire [16:0] mulnw_489;
wire [35:0] mul_678;
wire [15:0] mulnw_221;
wire [35:0] mul_410;
wire [17:0] add_599;
wire [15:0] slice_788;
wire [35:0] mul_142;
wire [40:0] subW_331;
wire [17:0] slice_520;
wire [17:0] add_709;
wire [17:0] slice_252;
wire [17:0] add_441;
wire [34:0] addW_630;
wire [50:0] addW_819;
wire [17:0] add_173;
wire [8:0] slice_362;
wire [71:0] subW_551;
wire [66:0] addW_740;
wire [8:0] slice_94;
wire [51:0] addW_283;
wire [16:0] slice_472;
wire [17:0] slice_661;
wire [196:0] addW_850;
wire [65:0] addW_204;
wire [17:0] slice_393;
wire [7:0] slice_582;
wire [7:0] slice_771;
wire [17:0] slice_125;
wire [41:0] subW_314;
wire [17:0] add_503;
wire [16:0] slice_692;
wire [27:0] mul_46;
wire [7:0] slice_235;
wire [16:0] slice_424;
wire [17:0] slice_613;
wire [15:0] mul_802;
wire [16:0] slice_156;
wire [31:0] mul_345;
wire [34:0] addW_534;
wire [25:0] lsl_723;
wire [25:0] lsl_455;
wire [17:0] slice_644;
wire [17:0] slice_833;
wire [25:0] lsl_187;
wire [15:0] slice_376;
wire [64:0] slice_565;
wire [16:0] mulnw_754;
wire [15:0] slice_108;
wire [63:0] slice_297;
wire [7:0] slice_486;
wire [27:0] mul_675;
wire [16:0] mulnw_218;
wire [27:0] mul_407;
wire [16:0] mulnw_596;
wire [16:0] slice_785;
wire [27:0] mul_139;
wire [19:0] addW_328;
wire [17:0] slice_517;
wire [15:0] mulnw_706;
wire [31:0] slice_60;
wire [13:0] slice_249;
wire [15:0] mulnw_438;
wire [98:0] concat_627;
wire [26:0] add_816;
wire [15:0] mulnw_170;
wire [26:0] add_359;
wire [17:0] slice_548;
wire [195:0] concat_737;
wire [26:0] add_91;
wire [39:0] mul_280;
wire [194:0] concat_469;
wire [17:0] slice_658;
wire [133:0] concat_847;
wire [194:0] concat_201;
wire [17:0] slice_390;
wire [7:0] slice_579;
wire [32:0] lsl_768;
wire [17:0] slice_122;
wire [19:0] addW_311;
wire [16:0] mulnw_500;
wire [31:0] slice_689;
wire [13:0] slice_43;
wire [32:0] lsl_232;
wire [31:0] slice_421;
wire [31:0] slice_610;
wire [16:0] mulnw_799;
wire [31:0] slice_153;
wire [33:0] mul_342;
wire [98:0] concat_531;
wire [7:0] slice_720;
wire [31:0] mul_74;
wire [65:0] concat_263;
wire [7:0] slice_452;
wire [40:0] subW_641;
wire [17:0] slice_830;
wire [7:0] slice_184;
wire [33:0] add_373;
wire [49:0] concat_751;
wire [33:0] add_105;
wire [63:0] slice_294;
wire [7:0] slice_483;
wire [13:0] slice_672;
wire [17:0] slice_26;
wire [49:0] concat_215;
wire [13:0] slice_404;
wire [16:0] mulnw_593;
wire [32:0] slice_782;
wire [13:0] slice_136;
wire [35:0] mul_325;
wire [31:0] slice_514;
wire [16:0] mulnw_703;
wire [47:0] addW_57;
wire [31:0] slice_246;
wire [16:0] mulnw_435;
wire [17:0] slice_624;
wire [17:0] add_813;
wire [16:0] mulnw_167;
wire [17:0] add_356;
wire [40:0] subW_545;
wire [31:0] slice_734;
wire [17:0] add_88;
wire [49:0] concat_277;
wire [31:0] slice_466;
wire [31:0] slice_655;
wire [71:0] subW_844;
wire [31:0] slice_198;
wire [31:0] slice_387;
wire [15:0] slice_576;
wire [7:0] slice_765;
wire [31:0] slice_119;
wire [17:0] slice_308;
wire [16:0] mulnw_497;
wire [47:0] addW_686;
wire [17:0] slice_40;
wire [7:0] slice_229;
wire [47:0] addW_418;
wire [66:0] concat_607;
wire [7:0] slice_796;
wire [47:0] addW_150;
wire [16:0] slice_339;
wire [17:0] slice_528;
wire [32:0] lsl_717;
wire [41:0] subW_260;
wire [32:0] lsl_449;
wire [19:0] addW_638;
wire [34:0] addW_827;
wire [32:0] lsl_181;
wire [25:0] lsl_370;
wire [259:0] concat_559;
wire [15:0] slice_748;
wire [25:0] lsl_102;
wire [132:0] subW_291;
wire [15:0] slice_480;
wire [17:0] slice_669;
wire [27:0] mul_23;
wire [15:0] slice_212;
wire [17:0] slice_401;
wire [33:0] add_590;
wire [50:0] addW_779;
wire [17:0] slice_133;
wire [27:0] mul_322;
wire [66:0] concat_511;
wire [49:0] concat_700;
wire [39:0] mul_54;
wire [50:0] addW_243;
wire [49:0] concat_432;
wire [40:0] subW_621;
wire [16:0] mulnw_810;
wire [49:0] concat_164;
wire [15:0] mulnw_353;
wire [19:0] addW_542;
wire [67:0] subW_731;
wire [15:0] mulnw_85;
wire [17:0] slice_274;
wire [67:0] subW_463;
wire [31:0] slice_652;
wire [17:0] slice_841;
wire [67:0] subW_195;
wire [31:0] slice_384;
wire [15:0] slice_573;
wire [15:0] mul_762;
wire [31:0] slice_116;
wire [17:0] slice_305;
wire [33:0] add_494;
wire [39:0] mul_683;
wire [40:0] subW_37;
wire [15:0] mul_226;
wire [39:0] mul_415;
wire [34:0] addW_604;
wire [7:0] slice_793;
wire [39:0] mul_147;
wire [31:0] slice_336;
wire [40:0] subW_525;
wire [7:0] slice_714;
wire [33:0] addW_68;
wire [19:0] addW_257;
wire [7:0] slice_446;
wire [35:0] mul_635;
wire [7:0] slice_178;
wire [7:0] slice_367;
wire [133:0] subW_556;
wire [16:0] slice_745;
wire [7:0] slice_99;
wire [99:0] addW_288;
wire [15:0] slice_477;
wire [40:0] subW_666;
wire [388:0] addW_855;
wire [63:0] slice_20;
wire [16:0] slice_209;
wire [40:0] subW_398;
wire [25:0] lsl_587;
wire [26:0] add_776;
wire [40:0] subW_130;
wire [13:0] slice_319;
wire [34:0] addW_508;
wire [15:0] slice_697;
wire [45:0] concat_51;
wire [26:0] add_240;
wire [15:0] slice_429;
wire [19:0] addW_618;
wire [16:0] mulnw_807;
wire [15:0] slice_161;
wire [16:0] mulnw_350;
wire [35:0] mul_539;
wire [50:0] addW_728;
wire [32:0] lsl_82;
wire [15:0] slice_271;
wire [50:0] addW_460;
wire [31:0] slice_649;
wire [40:0] subW_838;
wire [50:0] addW_192;
wire [31:0] slice_381;
wire [32:0] slice_570;
wire [16:0] mulnw_759;
wire [31:0] slice_113;
wire [31:0] slice_302;
wire [25:0] lsl_491;
wire [45:0] concat_680;
wire [19:0] addW_34;
wire [16:0] mulnw_223;
wire [45:0] concat_412;
wire [15:0] mul_601;
wire [15:0] slice_790;
wire [45:0] concat_144;
wire [47:0] addW_333;
wire [19:0] addW_522;
wire [15:0] mul_711;
wire [33:0] addW_65;
wire [17:0] slice_254;
wire [15:0] mul_443;
wire [31:0] mul_632;
wire [66:0] concat_821;
wire [15:0] mul_175;
wire [32:0] lsl_364;
wire [31:0] slice_553;
wire [16:0] slice_742;
wire [32:0] lsl_96;
wire [69:0] concat_285;
wire [32:0] slice_474;
wire [19:0] addW_663;
wire [260:0] concat_852;
wire [13:0] slice_17;
wire [16:0] slice_206;
wire [19:0] addW_395;
wire [7:0] slice_584;
wire [17:0] add_773;
wire [19:0] addW_127;
wire [17:0] slice_316;
wire [15:0] mul_505;
wire [16:0] slice_694;
wire [17:0] slice_48;
wire [17:0] add_237;
wire [16:0] slice_426;
wire [35:0] mul_615;
wire [33:0] add_804;
wire [16:0] slice_158;
wire [49:0] concat_347;
wire [31:0] mul_536;
wire [26:0] add_725;
wire [8:0] slice_79;
wire [34:0] addW_268;
wire [26:0] add_457;
wire [70:0] subW_646;
wire [19:0] addW_835;
assign add_189 = lsl_187 + mul_188;
assign subW_378 = concat_377 - concat_317;
assign slice_567 = slice_566[32:16];
assign slice_756 = slice_742[7:0];
assign subW_110 = concat_109 - concat_41;
assign slice_299 = slice_298[31:18];
assign slice_488 = slice_478[7:0];
assign slice_677 = slice_673[17:0];
assign concat_31 = {mul_23,slice_30};
assign slice_220 = slice_206[7:0];
assign slice_409 = slice_405[17:0];
assign mulnw_598 = slice_591 * slice_597;
assign slice_787 = slice_782[15:0];
assign slice_141 = slice_137[17:0];
assign mul_330 = addW_328 * addW_329;
assign mul_519 = slice_517 * slice_518;
assign mulnw_708 = slice_701 * slice_707;
assign slice_251 = slice_246[17:0];
assign mulnw_440 = slice_433 * slice_439;
assign slice_629 = addW_628[33:18];
assign addW_818 = add_804 + add_817;
assign mulnw_172 = slice_165 * slice_171;
assign slice_361 = slice_343[15:8];
assign subW_550 = concat_549 - concat_511;
assign slice_93 = slice_72[15:8];
assign subW_282 = subW_281 - mul_275;
assign slice_471 = addW_470[64:32];
assign mul_660 = slice_658 * slice_659;
assign subW_849 = subW_848 - concat_735;
assign slice_14 = slice_11[63:32];
assign mul_392 = slice_390 * slice_391;
assign lsl_581 = mulnw_580 << 16;
assign mulnw_770 = slice_769 * slice_766;
assign mul_124 = slice_122 * slice_123;
assign subW_313 = mul_312 - mul_304;
assign mulnw_502 = slice_495 * slice_501;
assign addW_691 = slice_671 + slice_652;
assign slice_45 = slice_44[31:18];
assign mulnw_234 = slice_233 * slice_230;
assign addW_423 = slice_403 + slice_384;
assign mul_612 = slice_609 * slice_611;
assign lsl_801 = add_800 << 8;
assign addW_155 = slice_135 + slice_116;
assign slice_344 = addW_340[15:0];
assign slice_533 = addW_532[33:18];
assign add_722 = mulnw_719 + mulnw_721;
assign concat_76 = {mul_70,slice_75};
assign concat_265 = {concat_245,slice_264};
assign add_454 = mulnw_451 + mulnw_453;
assign addW_643 = concat_637 + subW_642;
assign mul_832 = slice_830 * slice_831;
assign add_186 = mulnw_183 + mulnw_185;
assign addW_375 = concat_347 + addW_374;
assign addW_564 = slice_296 + slice_8;
assign slice_753 = slice_748[15:8];
assign addW_107 = concat_76 + addW_106;
assign slice_296 = IN1[127:0];
assign lsl_485 = mulnw_484 << 16;
assign slice_674 = slice_673[31:18];
assign mul_28 = slice_26 * slice_27;
assign slice_217 = slice_212[15:8];
assign slice_406 = slice_405[31:18];
assign slice_595 = slice_573[7:0];
assign slice_784 = addW_743[32:0];
assign slice_138 = slice_137[31:18];
assign concat_327 = {mul_322,slice_326};
assign mul_516 = slice_513 * slice_515;
assign slice_705 = slice_692[7:0];
assign concat_59 = {addW_57,slice_58};
assign slice_248 = addW_207[31:0];
assign slice_437 = slice_424[7:0];
assign slice_626 = concat_625[63:32];
assign mul_815 = slice_809 * slice_811;
assign slice_169 = slice_156[7:0];
assign mul_358 = slice_352 * slice_354;
assign addW_547 = concat_541 + subW_546;
assign slice_736 = concat_735[127:64];
assign mul_90 = slice_84 * slice_86;
assign addW_279 = slice_274 + slice_271;
assign slice_468 = concat_467[127:64];
assign mul_657 = slice_653 * slice_656;
assign slice_846 = concat_821[32:0];
assign slice_11 = slice_8[127:64];
assign slice_200 = concat_199[127:64];
assign mul_389 = slice_385 * slice_388;
assign slice_578 = slice_567[16:8];
assign mulnw_767 = slice_765 * slice_766;
assign mul_121 = slice_117 * slice_120;
assign addW_310 = slice_305 + slice_299;
assign slice_499 = slice_477[7:0];
assign concat_688 = {addW_686,slice_687};
assign slice_42 = slice_11[31:0];
assign mulnw_231 = slice_229 * slice_230;
assign concat_420 = {addW_418,slice_419};
assign slice_609 = slice_608[31:18];
assign slice_798 = slice_788[7:0];
assign concat_152 = {addW_150,slice_151};
assign slice_341 = addW_340[32:16];
assign slice_530 = concat_529[63:32];
assign mulnw_719 = slice_718 * slice_715;
assign slice_73 = addW_68[15:0];
assign slice_262 = mul_253[17:0];
assign mulnw_451 = slice_450 * slice_447;
assign mul_640 = addW_638 * addW_639;
assign mul_829 = slice_826 * slice_828;
assign mulnw_183 = slice_182 * slice_179;
assign add_372 = lsl_370 + mul_371;
assign concat_561 = {concat_295,slice_560};
assign slice_750 = mul_749[31:16];
assign add_104 = lsl_102 + mul_103;
assign addW_293 = concat_201 + subW_292;
assign slice_482 = slice_472[16:8];
assign slice_671 = slice_651[31:0];
assign slice_214 = mul_213[31:16];
assign slice_403 = slice_383[31:0];
assign slice_592 = slice_571[16:8];
assign concat_781 = {addW_779,slice_780};
assign slice_135 = slice_115[31:0];
assign slice_324 = slice_320[17:0];
assign slice_513 = slice_512[31:18];
assign slice_702 = slice_697[15:8];
assign subW_56 = subW_55 - mul_49;
assign concat_245 = {addW_243,slice_244};
assign slice_434 = slice_429[15:8];
assign addW_623 = concat_617 + subW_622;
assign mulnw_812 = slice_805 * slice_811;
assign slice_166 = slice_161[15:8];
assign mulnw_355 = slice_348 * slice_354;
assign mul_544 = addW_542 * addW_543;
assign addW_733 = concat_690 + subW_732;
assign mulnw_87 = slice_79 * slice_86;
assign slice_276 = mul_275[35:18];
assign addW_465 = concat_422 + subW_464;
assign slice_654 = addW_568[63:0];
assign subW_843 = concat_842 - concat_781;
assign slice_8 = IN1[255:128];
assign addW_197 = concat_154 + subW_196;
assign slice_386 = slice_300[63:0];
assign mul_575 = slice_573 * slice_574;
assign add_764 = lsl_755 + add_763;
assign slice_118 = slice_19[63:0];
assign mul_307 = slice_305 * slice_306;
assign slice_496 = slice_475[16:8];
assign subW_685 = subW_684 - mul_678;
assign addW_39 = concat_31 + subW_38;
assign add_228 = lsl_219 + add_227;
assign subW_417 = subW_416 - mul_410;
assign slice_606 = mul_575[15:0];
assign lsl_795 = mulnw_794 << 16;
assign subW_149 = subW_148 - mul_142;
assign addW_338 = slice_318 + slice_298;
assign addW_527 = concat_521 + subW_526;
assign mulnw_716 = slice_714 * slice_715;
assign mul_70 = slice_67 * slice_69;
assign subW_259 = mul_258 - mul_250;
assign mulnw_448 = slice_446 * slice_447;
assign concat_637 = {mul_632,slice_636};
assign slice_826 = addW_825[33:18];
assign mulnw_180 = slice_178 * slice_179;
assign add_369 = mulnw_366 + mulnw_368;
assign slice_558 = concat_467[63:0];
assign slice_747 = slice_741[15:0];
assign add_101 = mulnw_98 + mulnw_100;
assign concat_290 = {addW_288,slice_289};
assign mul_479 = slice_477 * slice_478;
assign addW_668 = concat_662 + subW_667;
assign concat_857 = {addW_855,slice_856};
assign slice_22 = slice_21[31:18];
assign slice_211 = slice_205[15:0];
assign addW_400 = concat_394 + subW_399;
assign add_589 = lsl_587 + mul_588;
assign addW_778 = add_764 + add_777;
assign addW_132 = concat_126 + subW_131;
assign slice_321 = slice_320[31:18];
assign slice_510 = mul_479[15:0];
assign slice_699 = mul_698[31:16];
assign addW_53 = slice_48 + slice_45;
assign addW_242 = add_228 + add_241;
assign slice_431 = mul_430[31:16];
assign mul_620 = addW_618 * addW_619;
assign slice_809 = slice_787[7:0];
assign slice_163 = mul_162[31:16];
assign slice_352 = slice_339[7:0];
assign concat_541 = {mul_536,slice_540};
assign concat_730 = {addW_728,slice_729};
assign slice_84 = slice_67[7:0];
assign slice_273 = addW_268[17:0];
assign concat_462 = {addW_460,slice_461};
assign slice_651 = addW_564[63:0];
assign addW_840 = concat_834 + subW_839;
assign concat_194 = {addW_192,slice_193};
assign slice_383 = slice_296[63:0];
assign mul_572 = slice_567 * slice_571;
assign lsl_761 = add_760 << 8;
assign slice_115 = slice_8[63:0];
assign mul_304 = slice_299 * slice_303;
assign add_493 = lsl_491 + mul_492;
assign addW_682 = slice_677 + slice_674;
assign mul_36 = addW_34 * addW_35;
assign lsl_225 = add_224 << 8;
assign addW_414 = slice_409 + slice_406;
assign add_603 = lsl_594 + add_602;
assign slice_792 = slice_783[16:8];
assign addW_146 = slice_141 + slice_138;
assign concat_335 = {addW_333,slice_334};
assign mul_524 = addW_522 * addW_523;
assign add_713 = lsl_704 + add_712;
assign slice_67 = addW_65[32:16];
assign addW_256 = slice_251 + slice_247;
assign add_445 = lsl_436 + add_444;
assign slice_634 = addW_630[17:0];
assign concat_823 = {concat_781,slice_822};
assign add_177 = lsl_168 + add_176;
assign mulnw_366 = slice_365 * slice_362;
assign subW_555 = concat_554 - concat_382;
assign slice_744 = addW_743[65:33];
assign mulnw_98 = slice_97 * slice_94;
assign subW_287 = subW_286 - concat_263;
assign mul_476 = slice_472 * slice_475;
assign mul_665 = addW_663 * addW_664;
assign subW_854 = subW_853 - concat_559;
assign slice_19 = IN2[255:128];
assign slice_208 = addW_207[64:32];
assign mul_397 = addW_395 * addW_396;
assign add_586 = mulnw_583 + mulnw_585;
assign mul_775 = slice_769 * slice_771;
assign mul_129 = addW_127 * addW_128;
assign slice_318 = slice_297[31:0];
assign add_507 = lsl_498 + add_506;
assign slice_696 = addW_691[15:0];
assign slice_50 = mul_49[35:18];
assign mul_239 = slice_233 * slice_235;
assign slice_428 = addW_423[15:0];
assign concat_617 = {mul_612,slice_616};
assign slice_806 = slice_785[16:8];
assign slice_160 = addW_155[15:0];
assign slice_349 = slice_344[15:8];
assign slice_538 = addW_534[17:0];
assign addW_727 = add_713 + add_726;
assign mulnw_81 = slice_79 * slice_80;
assign addW_270 = slice_248 + slice_208;
assign addW_459 = add_445 + add_458;
assign addW_648 = concat_627 + subW_647;
assign mul_837 = addW_835 * addW_836;
assign addW_191 = add_177 + add_190;
assign addW_380 = concat_337 + subW_379;
assign slice_569 = addW_568[128:64];
assign slice_758 = slice_748[7:0];
assign addW_112 = concat_61 + subW_111;
assign slice_301 = slice_300[127:64];
assign add_490 = mulnw_487 + mulnw_489;
assign slice_679 = mul_678[35:18];
assign slice_222 = slice_212[7:0];
assign slice_411 = mul_410[35:18];
assign lsl_600 = add_599 << 8;
assign mul_789 = slice_787 * slice_788;
assign slice_143 = mul_142[35:18];
assign subW_332 = subW_331 - mul_325;
assign concat_521 = {mul_516,slice_520};
assign lsl_710 = add_709 << 8;
assign mul_253 = slice_251 * slice_252;
assign lsl_442 = add_441 << 8;
assign slice_631 = addW_630[33:18];
assign slice_820 = mul_789[15:0];
assign lsl_174 = add_173 << 8;
assign mulnw_363 = slice_361 * slice_362;
assign addW_552 = concat_531 + subW_551;
assign slice_741 = addW_740[65:33];
assign mulnw_95 = slice_93 * slice_94;
assign slice_284 = mul_275[17:0];
assign addW_473 = slice_386 + slice_301;
assign concat_662 = {mul_657,slice_661};
assign slice_851 = concat_735[63:0];
assign slice_205 = addW_204[64:32];
assign concat_394 = {mul_389,slice_393};
assign mulnw_583 = slice_582 * slice_579;
assign mulnw_772 = slice_765 * slice_771;
assign concat_126 = {mul_121,slice_125};
assign addW_315 = concat_309 + subW_314;
assign lsl_504 = add_503 << 8;
assign addW_693 = slice_673 + slice_655;
assign slice_47 = slice_42[17:0];
assign mulnw_236 = slice_229 * slice_235;
assign addW_425 = slice_405 + slice_387;
assign slice_614 = slice_610[17:0];
assign add_803 = lsl_801 + mul_802;
assign addW_157 = slice_137 + slice_119;
assign slice_346 = mul_345[31:16];
assign slice_535 = addW_534[33:18];
assign mul_724 = slice_718 * slice_720;
assign mul_456 = slice_450 * slice_452;
assign concat_645 = {addW_643,slice_644};
assign concat_834 = {mul_829,slice_833};
assign mul_188 = slice_182 * slice_184;
assign concat_377 = {addW_375,slice_376};
assign slice_566 = slice_565[64:32];
assign lsl_755 = mulnw_754 << 16;
assign concat_109 = {addW_107,slice_108};
assign slice_298 = slice_297[63:32];
assign mulnw_487 = slice_486 * slice_483;
assign slice_676 = slice_671[17:0];
assign slice_30 = mul_28[35:18];
assign lsl_219 = mulnw_218 << 16;
assign slice_408 = slice_403[17:0];
assign slice_597 = slice_571[7:0];
assign mul_786 = slice_783 * slice_785;
assign slice_140 = slice_135[17:0];
assign addW_329 = slice_324 + slice_321;
assign slice_518 = slice_514[17:0];
assign slice_707 = slice_697[7:0];
assign concat_61 = {concat_41,slice_60};
assign mul_250 = slice_247 * slice_249;
assign slice_439 = slice_429[7:0];
assign addW_628 = slice_608 + slice_566;
assign add_817 = lsl_808 + add_816;
assign slice_171 = slice_161[7:0];
assign add_360 = lsl_351 + add_359;
assign concat_549 = {addW_547,slice_548};
assign add_92 = lsl_82 + add_91;
assign subW_281 = mul_280 - mul_272;
assign addW_470 = slice_383 + slice_297;
assign slice_659 = slice_655[17:0];
assign subW_848 = concat_847 - concat_650;
assign slice_391 = slice_387[17:0];
assign mulnw_580 = slice_578 * slice_579;
assign slice_769 = slice_747[7:0];
assign slice_123 = slice_119[17:0];
assign mul_312 = addW_310 * addW_311;
assign slice_501 = slice_475[7:0];
assign concat_690 = {concat_670,slice_689};
assign slice_44 = slice_20[31:0];
assign slice_233 = slice_211[7:0];
assign concat_422 = {concat_402,slice_421};
assign slice_611 = slice_610[31:18];
assign add_800 = mulnw_797 + mulnw_799;
assign concat_154 = {concat_134,slice_153};
assign slice_343 = addW_338[15:0];
assign addW_532 = slice_512 + slice_471;
assign mulnw_721 = slice_714 * slice_720;
assign slice_75 = mul_74[31:16];
assign slice_264 = concat_263[63:32];
assign mulnw_453 = slice_446 * slice_452;
assign subW_642 = subW_641 - mul_635;
assign slice_831 = addW_827[17:0];
assign mulnw_185 = slice_178 * slice_184;
assign addW_374 = add_360 + add_373;
assign slice_752 = slice_742[16:8];
assign addW_106 = add_92 + add_105;
assign concat_295 = {addW_293,slice_294};
assign mulnw_484 = slice_482 * slice_483;
assign slice_673 = slice_654[31:0];
assign slice_27 = slice_21[17:0];
assign slice_216 = slice_206[16:8];
assign slice_405 = slice_386[31:0];
assign lsl_594 = mulnw_593 << 16;
assign slice_783 = slice_782[32:16];
assign slice_137 = slice_118[31:0];
assign slice_326 = mul_325[35:18];
assign slice_515 = slice_514[31:18];
assign lsl_704 = mulnw_703 << 16;
assign slice_58 = mul_49[17:0];
assign slice_247 = slice_246[31:18];
assign lsl_436 = mulnw_435 << 16;
assign concat_625 = {addW_623,slice_624};
assign lsl_814 = add_813 << 8;
assign lsl_168 = mulnw_167 << 16;
assign lsl_357 = add_356 << 8;
assign subW_546 = subW_545 - mul_539;
assign concat_735 = {addW_733,slice_734};
assign lsl_89 = add_88 << 8;
assign addW_278 = slice_273 + slice_269;
assign concat_467 = {addW_465,slice_466};
assign slice_656 = slice_655[31:18];
assign addW_845 = concat_823 + subW_844;
assign concat_199 = {addW_197,slice_198};
assign slice_388 = slice_387[31:18];
assign concat_577 = {mul_572,slice_576};
assign slice_766 = slice_745[16:8];
assign slice_120 = slice_119[31:18];
assign concat_309 = {mul_304,slice_308};
assign lsl_498 = mulnw_497 << 16;
assign slice_687 = mul_678[17:0];
assign concat_41 = {addW_39,slice_40};
assign slice_230 = slice_209[16:8];
assign slice_419 = mul_410[17:0];
assign slice_608 = slice_565[31:0];
assign mulnw_797 = slice_796 * slice_793;
assign slice_151 = mul_142[17:0];
assign addW_340 = slice_320 + slice_302;
assign concat_529 = {addW_527,slice_528};
assign slice_718 = slice_696[7:0];
assign slice_72 = addW_65[15:0];
assign addW_261 = concat_255 + subW_260;
assign slice_450 = slice_428[7:0];
assign addW_639 = slice_634 + slice_631;
assign slice_828 = addW_827[33:18];
assign slice_182 = slice_160[7:0];
assign mul_371 = slice_365 * slice_367;
assign slice_560 = concat_559[255:128];
assign mul_749 = slice_747 * slice_748;
assign mul_103 = slice_97 * slice_99;
assign subW_292 = subW_291 - concat_199;
assign concat_481 = {mul_476,slice_480};
assign concat_670 = {addW_668,slice_669};
assign mul_213 = slice_211 * slice_212;
assign concat_402 = {addW_400,slice_401};
assign slice_591 = slice_573[15:8];
assign slice_780 = mul_749[15:0];
assign concat_134 = {addW_132,slice_133};
assign slice_323 = slice_318[17:0];
assign slice_512 = addW_470[31:0];
assign slice_701 = slice_692[16:8];
assign subW_55 = mul_54 - mul_46;
assign slice_244 = mul_213[15:0];
assign slice_433 = slice_424[16:8];
assign subW_622 = subW_621 - mul_615;
assign slice_811 = slice_785[7:0];
assign slice_165 = slice_156[16:8];
assign slice_354 = slice_344[7:0];
assign addW_543 = slice_538 + slice_535;
assign subW_732 = subW_731 - concat_688;
assign slice_86 = slice_73[7:0];
assign mul_275 = slice_273 * slice_274;
assign subW_464 = subW_463 - concat_420;
assign slice_653 = slice_652[31:18];
assign concat_842 = {addW_840,slice_841};
assign subW_196 = subW_195 - concat_152;
assign slice_385 = slice_384[31:18];
assign slice_574 = slice_570[15:0];
assign add_763 = lsl_761 + mul_762;
assign slice_117 = slice_116[31:18];
assign slice_306 = slice_302[17:0];
assign slice_495 = slice_477[15:8];
assign subW_684 = mul_683 - mul_675;
assign subW_38 = subW_37 - mul_28;
assign add_227 = lsl_225 + mul_226;
assign subW_416 = mul_415 - mul_407;
assign addW_605 = concat_577 + addW_604;
assign mulnw_794 = slice_792 * slice_793;
assign subW_148 = mul_147 - mul_139;
assign concat_337 = {concat_317,slice_336};
assign subW_526 = subW_525 - mul_519;
assign slice_715 = slice_694[16:8];
assign slice_69 = addW_68[32:16];
assign mul_258 = addW_256 * addW_257;
assign slice_447 = slice_426[16:8];
assign slice_636 = mul_635[35:18];
assign addW_825 = slice_782 + slice_741;
assign slice_179 = slice_158[16:8];
assign mulnw_368 = slice_361 * slice_367;
assign addW_557 = concat_469 + subW_556;
assign mul_746 = slice_742 * slice_745;
assign mulnw_100 = slice_93 * slice_99;
assign slice_289 = concat_263[31:0];
assign slice_478 = slice_474[15:0];
assign subW_667 = subW_666 - mul_660;
assign slice_856 = concat_559[127:0];
assign slice_21 = slice_20[63:32];
assign mul_210 = slice_206 * slice_209;
assign subW_399 = subW_398 - mul_392;
assign mul_588 = slice_582 * slice_584;
assign add_777 = lsl_768 + add_776;
assign subW_131 = subW_130 - mul_124;
assign slice_320 = slice_301[31:0];
assign addW_509 = concat_481 + addW_508;
assign mul_698 = slice_696 * slice_697;
assign addW_52 = slice_47 + slice_43;
assign add_241 = lsl_232 + add_240;
assign mul_430 = slice_428 * slice_429;
assign addW_619 = slice_614 + slice_611;
assign lsl_808 = mulnw_807 << 16;
assign mul_162 = slice_160 * slice_161;
assign lsl_351 = mulnw_350 << 16;
assign slice_540 = mul_539[35:18];
assign slice_729 = mul_698[15:0];
assign mul_272 = slice_269 * slice_271;
assign slice_461 = mul_430[15:0];
assign concat_650 = {addW_648,slice_649};
assign subW_839 = subW_838 - mul_832;
assign slice_193 = mul_162[15:0];
assign concat_382 = {addW_380,slice_381};
assign slice_571 = slice_570[32:16];
assign add_760 = mulnw_757 + mulnw_759;
assign concat_114 = {addW_112,slice_113};
assign slice_303 = slice_302[31:18];
assign mul_492 = slice_486 * slice_488;
assign addW_681 = slice_676 + slice_672;
assign addW_35 = slice_27 + slice_22;
assign add_224 = mulnw_221 + mulnw_223;
assign addW_413 = slice_408 + slice_404;
assign add_602 = lsl_600 + mul_601;
assign concat_791 = {mul_786,slice_790};
assign addW_145 = slice_140 + slice_136;
assign slice_334 = mul_325[17:0];
assign addW_523 = slice_518 + slice_515;
assign add_712 = lsl_710 + mul_711;
assign concat_255 = {mul_250,slice_254};
assign add_444 = lsl_442 + mul_443;
assign slice_633 = addW_628[17:0];
assign slice_822 = concat_821[65:33];
assign add_176 = lsl_174 + mul_175;
assign slice_365 = slice_343[7:0];
assign concat_554 = {addW_552,slice_553};
assign addW_743 = slice_654 + slice_569;
assign slice_97 = slice_72[7:0];
assign subW_286 = concat_285 - concat_245;
assign slice_475 = slice_474[32:16];
assign addW_664 = slice_659 + slice_656;
assign subW_853 = concat_852 - concat_295;
assign addW_207 = slice_118 + slice_20;
assign addW_396 = slice_391 + slice_388;
assign mulnw_585 = slice_578 * slice_584;
assign lsl_774 = add_773 << 8;
assign addW_128 = slice_123 + slice_120;
assign concat_317 = {addW_315,slice_316};
assign add_506 = lsl_504 + mul_505;
assign mul_695 = slice_692 * slice_694;
assign mul_49 = slice_47 * slice_48;
assign lsl_238 = add_237 << 8;
assign mul_427 = slice_424 * slice_426;
assign slice_616 = mul_615[35:18];
assign slice_805 = slice_787[15:8];
assign mul_159 = slice_156 * slice_158;
assign slice_348 = slice_339[16:8];
assign slice_537 = addW_532[17:0];
assign add_726 = lsl_717 + add_725;
assign slice_80 = slice_73[15:8];
assign slice_269 = addW_268[33:18];
assign add_458 = lsl_449 + add_457;
assign subW_647 = subW_646 - concat_625;
assign addW_836 = slice_831 + slice_828;
assign add_190 = lsl_181 + add_189;
assign subW_379 = subW_378 - concat_335;
assign addW_568 = slice_300 + slice_19;
assign mulnw_757 = slice_756 * slice_753;
assign subW_111 = subW_110 - concat_59;
assign slice_300 = IN2[127:0];
assign mulnw_489 = slice_482 * slice_488;
assign mul_678 = slice_676 * slice_677;
assign mulnw_221 = slice_220 * slice_217;
assign mul_410 = slice_408 * slice_409;
assign add_599 = mulnw_596 + mulnw_598;
assign slice_788 = slice_784[15:0];
assign mul_142 = slice_140 * slice_141;
assign subW_331 = mul_330 - mul_322;
assign slice_520 = mul_519[35:18];
assign add_709 = mulnw_706 + mulnw_708;
assign slice_252 = slice_248[17:0];
assign add_441 = mulnw_438 + mulnw_440;
assign addW_630 = slice_610 + slice_570;
assign addW_819 = concat_791 + addW_818;
assign add_173 = mulnw_170 + mulnw_172;
assign slice_362 = slice_341[16:8];
assign subW_551 = subW_550 - concat_529;
assign addW_740 = slice_651 + slice_565;
assign slice_94 = slice_69[16:8];
assign addW_283 = concat_277 + subW_282;
assign slice_472 = slice_471[32:16];
assign slice_661 = mul_660[35:18];
assign addW_850 = concat_737 + subW_849;
assign addW_204 = slice_115 + slice_11;
assign slice_393 = mul_392[35:18];
assign slice_582 = slice_567[7:0];
assign slice_771 = slice_745[7:0];
assign slice_125 = mul_124[35:18];
assign subW_314 = subW_313 - mul_307;
assign add_503 = mulnw_500 + mulnw_502;
assign slice_692 = addW_691[32:16];
assign mul_46 = slice_43 * slice_45;
assign slice_235 = slice_209[7:0];
assign slice_424 = addW_423[32:16];
assign slice_613 = slice_608[17:0];
assign mul_802 = slice_796 * slice_798;
assign slice_156 = addW_155[32:16];
assign mul_345 = slice_343 * slice_344;
assign addW_534 = slice_514 + slice_474;
assign lsl_723 = add_722 << 8;
assign lsl_455 = add_454 << 8;
assign slice_644 = mul_635[17:0];
assign slice_833 = mul_832[35:18];
assign lsl_187 = add_186 << 8;
assign slice_376 = mul_345[15:0];
assign slice_565 = addW_564[128:64];
assign mulnw_754 = slice_752 * slice_753;
assign slice_108 = mul_74[15:0];
assign slice_297 = slice_296[127:64];
assign slice_486 = slice_472[7:0];
assign mul_675 = slice_672 * slice_674;
assign mulnw_218 = slice_216 * slice_217;
assign mul_407 = slice_404 * slice_406;
assign mulnw_596 = slice_595 * slice_592;
assign slice_785 = slice_784[32:16];
assign mul_139 = slice_136 * slice_138;
assign addW_328 = slice_323 + slice_319;
assign slice_517 = slice_512[17:0];
assign mulnw_706 = slice_705 * slice_702;
assign slice_60 = concat_59[63:32];
assign slice_249 = slice_248[31:18];
assign mulnw_438 = slice_437 * slice_434;
assign concat_627 = {concat_607,slice_626};
assign add_816 = lsl_814 + mul_815;
assign mulnw_170 = slice_169 * slice_166;
assign add_359 = lsl_357 + mul_358;
assign slice_548 = mul_539[17:0];
assign concat_737 = {concat_650,slice_736};
assign add_91 = lsl_89 + mul_90;
assign mul_280 = addW_278 * addW_279;
assign concat_469 = {concat_382,slice_468};
assign slice_658 = slice_652[17:0];
assign concat_847 = {addW_845,slice_846};
assign concat_201 = {concat_114,slice_200};
assign slice_390 = slice_384[17:0];
assign slice_579 = slice_574[15:8];
assign lsl_768 = mulnw_767 << 16;
assign slice_122 = slice_116[17:0];
assign addW_311 = slice_306 + slice_303;
assign mulnw_500 = slice_499 * slice_496;
assign slice_689 = concat_688[63:32];
assign slice_43 = slice_42[31:18];
assign lsl_232 = mulnw_231 << 16;
assign slice_421 = concat_420[63:32];
assign slice_610 = slice_569[31:0];
assign mulnw_799 = slice_792 * slice_798;
assign slice_153 = concat_152[63:32];
assign mul_342 = slice_339 * slice_341;
assign concat_531 = {concat_511,slice_530};
assign slice_720 = slice_694[7:0];
assign mul_74 = slice_72 * slice_73;
assign concat_263 = {addW_261,slice_262};
assign slice_452 = slice_426[7:0];
assign subW_641 = mul_640 - mul_632;
assign slice_830 = addW_825[17:0];
assign slice_184 = slice_158[7:0];
assign add_373 = lsl_364 + add_372;
assign concat_751 = {mul_746,slice_750};
assign add_105 = lsl_96 + add_104;
assign slice_294 = concat_199[63:0];
assign slice_483 = slice_478[15:8];
assign slice_672 = slice_671[31:18];
assign slice_26 = slice_14[17:0];
assign concat_215 = {mul_210,slice_214};
assign slice_404 = slice_403[31:18];
assign mulnw_593 = slice_591 * slice_592;
assign slice_782 = addW_740[32:0];
assign slice_136 = slice_135[31:18];
assign mul_325 = slice_323 * slice_324;
assign slice_514 = addW_473[31:0];
assign mulnw_703 = slice_701 * slice_702;
assign addW_57 = concat_51 + subW_56;
assign slice_246 = addW_204[31:0];
assign mulnw_435 = slice_433 * slice_434;
assign slice_624 = mul_615[17:0];
assign add_813 = mulnw_810 + mulnw_812;
assign mulnw_167 = slice_165 * slice_166;
assign add_356 = mulnw_353 + mulnw_355;
assign subW_545 = mul_544 - mul_536;
assign slice_734 = concat_688[31:0];
assign add_88 = mulnw_85 + mulnw_87;
assign concat_277 = {mul_272,slice_276};
assign slice_466 = concat_420[31:0];
assign slice_655 = slice_654[63:32];
assign subW_844 = subW_843 - concat_821;
assign slice_198 = concat_152[31:0];
assign slice_387 = slice_386[63:32];
assign slice_576 = mul_575[31:16];
assign slice_765 = slice_747[15:8];
assign slice_119 = slice_118[63:32];
assign slice_308 = mul_307[35:18];
assign mulnw_497 = slice_495 * slice_496;
assign addW_686 = concat_680 + subW_685;
assign slice_40 = mul_28[17:0];
assign slice_229 = slice_211[15:8];
assign addW_418 = concat_412 + subW_417;
assign concat_607 = {addW_605,slice_606};
assign slice_796 = slice_783[7:0];
assign addW_150 = concat_144 + subW_149;
assign slice_339 = addW_338[32:16];
assign slice_528 = mul_519[17:0];
assign lsl_717 = mulnw_716 << 16;
assign subW_260 = subW_259 - mul_253;
assign lsl_449 = mulnw_448 << 16;
assign addW_638 = slice_633 + slice_629;
assign addW_827 = slice_784 + slice_744;
assign lsl_181 = mulnw_180 << 16;
assign lsl_370 = add_369 << 8;
assign concat_559 = {addW_557,slice_558};
assign slice_748 = slice_744[15:0];
assign lsl_102 = add_101 << 8;
assign subW_291 = concat_290 - concat_114;
assign slice_480 = mul_479[31:16];
assign slice_669 = mul_660[17:0];
assign mul_23 = slice_17 * slice_22;
assign slice_212 = slice_208[15:0];
assign slice_401 = mul_392[17:0];
assign add_590 = lsl_581 + add_589;
assign addW_779 = concat_751 + addW_778;
assign slice_133 = mul_124[17:0];
assign mul_322 = slice_319 * slice_321;
assign concat_511 = {addW_509,slice_510};
assign concat_700 = {mul_695,slice_699};
assign mul_54 = addW_52 * addW_53;
assign addW_243 = concat_215 + addW_242;
assign concat_432 = {mul_427,slice_431};
assign subW_621 = mul_620 - mul_612;
assign mulnw_810 = slice_809 * slice_806;
assign concat_164 = {mul_159,slice_163};
assign mulnw_353 = slice_352 * slice_349;
assign addW_542 = slice_537 + slice_533;
assign subW_731 = concat_730 - concat_670;
assign mulnw_85 = slice_84 * slice_80;
assign slice_274 = addW_270[17:0];
assign subW_463 = concat_462 - concat_402;
assign slice_652 = slice_651[63:32];
assign slice_841 = mul_832[17:0];
assign subW_195 = concat_194 - concat_134;
assign slice_384 = slice_383[63:32];
assign slice_573 = slice_566[15:0];
assign mul_762 = slice_756 * slice_758;
assign slice_116 = slice_115[63:32];
assign slice_305 = slice_298[17:0];
assign add_494 = lsl_485 + add_493;
assign mul_683 = addW_681 * addW_682;
assign subW_37 = mul_36 - mul_23;
assign mul_226 = slice_220 * slice_222;
assign mul_415 = addW_413 * addW_414;
assign addW_604 = add_590 + add_603;
assign slice_793 = slice_788[15:8];
assign mul_147 = addW_145 * addW_146;
assign slice_336 = concat_335[63:32];
assign subW_525 = mul_524 - mul_516;
assign slice_714 = slice_696[15:8];
assign addW_68 = slice_44 + slice_21;
assign addW_257 = slice_252 + slice_249;
assign slice_446 = slice_428[15:8];
assign mul_635 = slice_633 * slice_634;
assign slice_178 = slice_160[15:8];
assign slice_367 = slice_341[7:0];
assign subW_556 = subW_555 - concat_467;
assign slice_745 = slice_744[32:16];
assign slice_99 = slice_69[7:0];
assign addW_288 = concat_265 + subW_287;
assign slice_477 = slice_471[15:0];
assign subW_666 = mul_665 - mul_657;
assign addW_855 = concat_561 + subW_854;
assign slice_20 = slice_19[127:64];
assign slice_209 = slice_208[32:16];
assign subW_398 = mul_397 - mul_389;
assign lsl_587 = add_586 << 8;
assign add_776 = lsl_774 + mul_775;
assign subW_130 = mul_129 - mul_121;
assign slice_319 = slice_318[31:18];
assign addW_508 = add_494 + add_507;
assign slice_697 = addW_693[15:0];
assign concat_51 = {mul_46,slice_50};
assign add_240 = lsl_238 + mul_239;
assign slice_429 = addW_425[15:0];
assign addW_618 = slice_613 + slice_609;
assign mulnw_807 = slice_805 * slice_806;
assign slice_161 = addW_157[15:0];
assign mulnw_350 = slice_348 * slice_349;
assign mul_539 = slice_537 * slice_538;
assign addW_728 = concat_700 + addW_727;
assign lsl_82 = mulnw_81 << 16;
assign slice_271 = addW_270[33:18];
assign addW_460 = concat_432 + addW_459;
assign slice_649 = concat_625[31:0];
assign subW_838 = mul_837 - mul_829;
assign addW_192 = concat_164 + addW_191;
assign slice_381 = concat_335[31:0];
assign slice_570 = slice_569[64:32];
assign mulnw_759 = slice_752 * slice_758;
assign slice_113 = concat_59[31:0];
assign slice_302 = slice_301[63:32];
assign lsl_491 = add_490 << 8;
assign concat_680 = {mul_675,slice_679};
assign addW_34 = slice_26 + slice_17;
assign mulnw_223 = slice_216 * slice_222;
assign concat_412 = {mul_407,slice_411};
assign mul_601 = slice_595 * slice_597;
assign slice_790 = mul_789[31:16];
assign concat_144 = {mul_139,slice_143};
assign addW_333 = concat_327 + subW_332;
assign addW_522 = slice_517 + slice_513;
assign mul_711 = slice_705 * slice_707;
assign addW_65 = slice_42 + slice_14;
assign slice_254 = mul_253[35:18];
assign mul_443 = slice_437 * slice_439;
assign mul_632 = slice_629 * slice_631;
assign concat_821 = {addW_819,slice_820};
assign mul_175 = slice_169 * slice_171;
assign lsl_364 = mulnw_363 << 16;
assign slice_553 = concat_529[31:0];
assign slice_742 = slice_741[32:16];
assign lsl_96 = mulnw_95 << 16;
assign concat_285 = {addW_283,slice_284};
assign slice_474 = addW_473[64:32];
assign addW_663 = slice_658 + slice_653;
assign concat_852 = {addW_850,slice_851};
assign slice_17 = slice_14[31:18];
assign slice_206 = slice_205[32:16];
assign addW_395 = slice_390 + slice_385;
assign slice_584 = slice_574[7:0];
assign add_773 = mulnw_770 + mulnw_772;
assign addW_127 = slice_122 + slice_117;
assign slice_316 = mul_307[17:0];
assign mul_505 = slice_499 * slice_501;
assign slice_694 = addW_693[32:16];
assign slice_48 = slice_44[17:0];
assign add_237 = mulnw_234 + mulnw_236;
assign slice_426 = addW_425[32:16];
assign mul_615 = slice_613 * slice_614;
assign add_804 = lsl_795 + add_803;
assign slice_158 = addW_157[32:16];
assign concat_347 = {mul_342,slice_346};
assign mul_536 = slice_533 * slice_535;
assign add_725 = lsl_723 + mul_724;
assign slice_79 = slice_67[16:8];
assign addW_268 = slice_246 + slice_205;
assign add_457 = lsl_455 + mul_456;
assign subW_646 = concat_645 - concat_607;
assign addW_835 = slice_830 + slice_826;
assign OUTPUT = concat_857;
    endmodule