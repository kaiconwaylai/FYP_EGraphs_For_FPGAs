//Alpha = 0.003. Cost: LUTs = 4644. DSPs = 0.  

`timescale 1ns / 1ps
    module mult(
        input[225:0] IN1,
        input[225:0] IN2,
        output[451:0] OUTPUT
    );
wire [5:0] slice_189;
wire [11:0] addW_378;
wire [13:0] slice_567;
wire [45:0] addW_756;
wire [19:0] addW_945;
wire [13:0] slice_1134;
wire [4:0] slice_1323;
wire [25:0] concat_1512;
wire [15:0] lsl_1701;
wire [13:0] mul_1890;
wire [41:0] subW_251;
wire [6:0] slice_440;
wire [17:0] slice_629;
wire [18:0] lsl_818;
wire [4:0] slice_1007;
wire [13:0] mul_1196;
wire [20:0] concat_1385;
wire [88:0] addW_1574;
wire [8:0] mulnw_1763;
wire [4:0] slice_1952;
wire [9:0] mul_124;
wire [8:0] mulnw_313;
wire [22:0] concat_502;
wire [118:0] concat_691;
wire [8:0] slice_880;
wire [8:0] slice_1069;
wire [45:0] addW_1258;
wire [4:0] slice_1447;
wire [59:0] concat_1636;
wire [13:0] mul_1825;
wire [5:0] slice_186;
wire [14:0] concat_375;
wire [23:0] addW_564;
wire [23:0] add_753;
wire [35:0] mul_942;
wire [29:0] add_1131;
wire [3:0] slice_1320;
wire [13:0] addW_1509;
wire [9:0] mulnw_1698;
wire [6:0] slice_1887;
wire [31:0] addW_248;
wire [6:0] slice_437;
wire [5:0] slice_626;
wire [19:0] add_815;
wire [4:0] slice_1004;
wire [13:0] mulnw_1193;
wire [6:0] slice_1382;
wire [62:0] concat_1571;
wire [8:0] slice_1760;
wire [4:0] slice_1949;
wire [19:0] addW_121;
wire [3:0] slice_310;
wire [6:0] slice_499;
wire [64:0] subW_688;
wire [4:0] slice_877;
wire [19:0] add_1066;
wire [23:0] add_1255;
wire [4:0] slice_1444;
wire [30:0] addW_1633;
wire [6:0] slice_1822;
wire [112:0] slice_2011;
wire [11:0] slice_183;
wire [4:0] slice_372;
wire [14:0] mul4_561;
wire [15:0] add_750;
wire [21:0] concat_939;
wire [22:0] lsl_1128;
wire [9:0] mul_1317;
wire [17:0] concat_1506;
wire [8:0] mulnw_1695;
wire [6:0] slice_1884;
wire [22:0] addW_56;
wire [16:0] add_245;
wire [14:0] mul4_434;
wire [11:0] mul_623;
wire [15:0] lsl_812;
wire [4:0] slice_1001;
wire [14:0] mulnw_1190;
wire [6:0] slice_1379;
wire [42:0] subW_1568;
wire [8:0] slice_1757;
wire [4:0] slice_1946;
wire [19:0] addW_118;
wire [17:0] mul_307;
wire [7:0] slice_496;
wire [17:0] slice_685;
wire [9:0] mul_874;
wire [15:0] lsl_1063;
wire [15:0] add_1252;
wire [4:0] slice_1441;
wire [13:0] mul_1630;
wire [6:0] slice_1819;
wire [232:0] subW_2008;
wire [11:0] slice_180;
wire [4:0] slice_369;
wire [13:0] mul_558;
wire [28:0] lsl_747;
wire [11:0] addW_936;
wire [14:0] mulnw_1125;
wire [9:0] mulnw_1314;
wire [5:0] slice_1503;
wire [16:0] add_1692;
wire [13:0] slice_1881;
wire [13:0] mul_53;
wire [10:0] add_242;
wire [6:0] slice_431;
wire [5:0] slice_620;
wire [4:0] slice_809;
wire [58:0] concat_998;
wire [13:0] mul_1187;
wire [13:0] slice_1376;
wire [8:0] slice_1565;
wire [16:0] addW_1754;
wire [43:0] concat_1943;
wire [39:0] concat_115;
wire [21:0] concat_304;
wire [58:0] addW_493;
wire [41:0] subW_682;
wire [4:0] slice_871;
wire [9:0] mulnw_1060;
wire [28:0] lsl_1249;
wire [39:0] concat_1438;
wire [13:0] mulnw_1627;
wire [14:0] mul4_1816;
wire [174:0] addW_2005;
wire [4:0] slice_366;
wire [15:0] mul_555;
wire [23:0] add_744;
wire [14:0] concat_933;
wire [29:0] add_1122;
wire [18:0] lsl_1311;
wire [5:0] slice_1500;
wire [10:0] add_1689;
wire [30:0] concat_1878;
wire [6:0] slice_50;
wire [4:0] slice_239;
wire [6:0] slice_428;
wire [5:0] slice_617;
wire [8:0] mulnw_806;
wire [42:0] subW_995;
wire [14:0] mulnw_1184;
wire [23:0] addW_1373;
wire [19:0] add_1562;
wire [9:0] mul_1751;
wire [17:0] slice_1940;
wire [35:0] mul_112;
wire [11:0] addW_301;
wire [28:0] slice_490;
wire [31:0] addW_679;
wire [4:0] slice_868;
wire [8:0] mulnw_1057;
wire [23:0] add_1246;
wire [17:0] slice_1435;
wire [14:0] mulnw_1624;
wire [6:0] slice_1813;
wire [118:0] concat_2002;
wire [39:0] concat_363;
wire [28:0] slice_552;
wire [15:0] add_741;
wire [4:0] slice_930;
wire [22:0] lsl_1119;
wire [30:0] concat_1308;
wire [5:0] slice_1497;
wire [8:0] mulnw_1686;
wire [16:0] addW_1875;
wire [6:0] slice_47;
wire [3:0] slice_236;
wire [14:0] slice_425;
wire [11:0] slice_614;
wire [8:0] slice_803;
wire [8:0] slice_992;
wire [14:0] mulnw_1181;
wire [14:0] mul4_1370;
wire [15:0] lsl_1559;
wire [9:0] mul_1748;
wire [5:0] slice_1937;
wire [14:0] concat_298;
wire [16:0] add_676;
wire [9:0] slice_865;
wire [16:0] add_1054;
wire [15:0] add_1243;
wire [4:0] slice_1432;
wire [13:0] mul_1621;
wire [6:0] slice_1810;
wire [64:0] subW_1999;
wire [40:0] addW_171;
wire [17:0] slice_360;
wire [28:0] slice_549;
wire [28:0] lsl_738;
wire [4:0] slice_927;
wire [13:0] mulnw_1116;
wire [8:0] slice_1305;
wire [87:0] concat_1494;
wire [3:0] slice_1683;
wire [22:0] concat_1872;
wire [13:0] slice_44;
wire [9:0] mul_233;
wire [14:0] slice_422;
wire [11:0] slice_611;
wire [8:0] slice_800;
wire [19:0] add_989;
wire [29:0] concat_1178;
wire [13:0] mul_1367;
wire [9:0] mulnw_1556;
wire [9:0] mul_1745;
wire [11:0] mul_1934;
wire [16:0] addW_106;
wire [4:0] slice_295;
wire [10:0] add_673;
wire [9:0] slice_862;
wire [10:0] add_1051;
wire [28:0] lsl_1240;
wire [9:0] mul_1429;
wire [14:0] mulnw_1618;
wire [14:0] slice_1807;
wire [17:0] slice_1996;
wire [40:0] concat_168;
wire [4:0] slice_357;
wire [45:0] addW_546;
wire [13:0] slice_735;
wire [55:0] slice_924;
wire [44:0] concat_1113;
wire [4:0] slice_1302;
wire [17:0] slice_1491;
wire [17:0] mul_1680;
wire [6:0] slice_1869;
wire [9:0] mulnw_230;
wire [86:0] concat_419;
wire [88:0] concat_608;
wire [16:0] addW_797;
wire [15:0] lsl_986;
wire [15:0] addW_1175;
wire [15:0] mul_1364;
wire [8:0] mulnw_1553;
wire [19:0] addW_1742;
wire [5:0] slice_1931;
wire [9:0] mul_103;
wire [4:0] slice_292;
wire [87:0] addW_481;
wire [4:0] slice_670;
wire [17:0] slice_859;
wire [8:0] mulnw_1048;
wire [13:0] slice_1237;
wire [4:0] slice_1426;
wire [14:0] mulnw_1615;
wire [7:0] slice_1804;
wire [41:0] subW_1993;
wire [20:0] addW_165;
wire [9:0] mul_354;
wire [23:0] add_543;
wire [22:0] addW_732;
wire [27:0] slice_921;
wire [6:0] slice_1110;
wire [9:0] mul_1299;
wire [41:0] subW_1488;
wire [21:0] concat_1677;
wire [7:0] slice_1866;
wire [23:0] addW_38;
wire [18:0] lsl_227;
wire [17:0] slice_416;
wire [13:0] slice_605;
wire [9:0] mul_794;
wire [9:0] mulnw_983;
wire [20:0] concat_1172;
wire [28:0] slice_1361;
wire [16:0] add_1550;
wire [19:0] addW_1739;
wire [5:0] slice_1928;
wire [4:0] slice_100;
wire [4:0] slice_289;
wire [59:0] concat_478;
wire [3:0] slice_667;
wire [17:0] slice_856;
wire [3:0] slice_1045;
wire [22:0] addW_1234;
wire [4:0] slice_1423;
wire [29:0] concat_1612;
wire [58:0] addW_1801;
wire [31:0] addW_1990;
wire [9:0] mul_162;
wire [4:0] slice_351;
wire [15:0] add_540;
wire [13:0] mul_729;
wire [27:0] slice_918;
wire [13:0] mul_1107;
wire [4:0] slice_1296;
wire [31:0] addW_1485;
wire [11:0] addW_1674;
wire [7:0] slice_1863;
wire [14:0] mul4_35;
wire [30:0] concat_224;
wire [41:0] subW_413;
wire [29:0] add_602;
wire [9:0] mul_791;
wire [8:0] mulnw_980;
wire [6:0] slice_1169;
wire [7:0] slice_1358;
wire [10:0] add_1547;
wire [35:0] mul_1736;
wire [11:0] slice_1925;
wire [4:0] slice_97;
wire [39:0] concat_286;
wire [30:0] addW_475;
wire [9:0] mul_664;
wire [19:0] addW_853;
wire [17:0] mul_1042;
wire [13:0] mul_1231;
wire [9:0] slice_1420;
wire [15:0] addW_1609;
wire [56:0] slice_1798;
wire [16:0] add_1987;
wire [8:0] mulnw_159;
wire [4:0] slice_348;
wire [28:0] lsl_537;
wire [13:0] mul_726;
wire [63:0] subW_915;
wire [6:0] slice_1104;
wire [4:0] slice_1293;
wire [16:0] add_1482;
wire [14:0] concat_1671;
wire [59:0] concat_1860;
wire [6:0] slice_32;
wire [8:0] slice_221;
wire [31:0] addW_410;
wire [22:0] lsl_599;
wire [9:0] mul_788;
wire [16:0] add_977;
wire [6:0] slice_1166;
wire [56:0] slice_1355;
wire [8:0] mulnw_1544;
wire [25:0] concat_1733;
wire [11:0] slice_1922;
wire [4:0] slice_94;
wire [17:0] slice_283;
wire [13:0] mul_472;
wire [9:0] mulnw_661;
wire [11:0] mul_850;
wire [21:0] concat_1039;
wire [13:0] mul_1228;
wire [9:0] slice_1417;
wire [20:0] concat_1606;
wire [88:0] addW_1795;
wire [10:0] add_1984;
wire [18:0] lsl_156;
wire [9:0] slice_345;
wire [23:0] add_534;
wire [13:0] mul_723;
wire [44:0] addW_912;
wire [6:0] slice_1101;
wire [9:0] slice_1290;
wire [10:0] add_1479;
wire [4:0] slice_1668;
wire [30:0] addW_1857;
wire [6:0] slice_29;
wire [4:0] slice_218;
wire [16:0] add_407;
wire [14:0] mulnw_596;
wire [19:0] addW_785;
wire [10:0] add_974;
wire [13:0] slice_1163;
wire [3:0] slice_1541;
wire [13:0] addW_1730;
wire [28:0] slice_1919;
wire [4:0] slice_91;
wire [4:0] slice_280;
wire [13:0] mulnw_469;
wire [18:0] lsl_658;
wire [11:0] mul_847;
wire [11:0] addW_1036;
wire [13:0] mul_1225;
wire [13:0] slice_1414;
wire [6:0] slice_1603;
wire [62:0] concat_1792;
wire [4:0] slice_1981;
wire [19:0] add_153;
wire [9:0] slice_342;
wire [15:0] add_531;
wire [6:0] slice_720;
wire [40:0] concat_909;
wire [13:0] slice_1098;
wire [9:0] slice_1287;
wire [4:0] slice_1476;
wire [4:0] slice_1665;
wire [13:0] mul_1854;
wire [9:0] mul_215;
wire [10:0] add_404;
wire [29:0] add_593;
wire [19:0] addW_782;
wire [8:0] mulnw_971;
wire [23:0] addW_1160;
wire [229:0] concat_1349;
wire [17:0] mul_1538;
wire [17:0] concat_1727;
wire [45:0] addW_1916;
wire [9:0] mul_277;
wire [14:0] mulnw_466;
wire [30:0] concat_655;
wire [11:0] mul_844;
wire [14:0] concat_1033;
wire [6:0] slice_1222;
wire [29:0] add_1411;
wire [6:0] slice_1600;
wire [42:0] subW_1789;
wire [3:0] slice_1978;
wire [15:0] lsl_150;
wire [17:0] slice_339;
wire [28:0] lsl_528;
wire [6:0] slice_717;
wire [20:0] addW_906;
wire [30:0] concat_1095;
wire [17:0] slice_1284;
wire [3:0] slice_1473;
wire [4:0] slice_1662;
wire [13:0] mulnw_1851;
wire [14:0] slice_23;
wire [4:0] slice_212;
wire [4:0] slice_401;
wire [22:0] lsl_590;
wire [35:0] mul_779;
wire [3:0] slice_968;
wire [14:0] mul4_1157;
wire [120:0] subW_1346;
wire [21:0] concat_1535;
wire [5:0] slice_1724;
wire [23:0] add_1913;
wire [4:0] slice_274;
wire [13:0] mul_463;
wire [8:0] slice_652;
wire [30:0] addW_841;
wire [4:0] slice_1030;
wire [6:0] slice_1219;
wire [22:0] lsl_1408;
wire [13:0] slice_1597;
wire [8:0] slice_1786;
wire [9:0] mul_1975;
wire [4:0] slice_147;
wire [41:0] subW_336;
wire [13:0] slice_525;
wire [14:0] mul4_714;
wire [9:0] mul_903;
wire [16:0] addW_1092;
wire [17:0] slice_1281;
wire [9:0] mul_1470;
wire [39:0] concat_1659;
wire [14:0] mulnw_1848;
wire [112:0] slice_20;
wire [4:0] slice_209;
wire [3:0] slice_398;
wire [13:0] mulnw_587;
wire [21:0] concat_776;
wire [17:0] mul_965;
wire [13:0] mul_1154;
wire [28:0] slice_1343;
wire [11:0] addW_1532;
wire [5:0] slice_1721;
wire [15:0] add_1910;
wire [45:0] addW_82;
wire [4:0] slice_271;
wire [14:0] mulnw_460;
wire [4:0] slice_649;
wire [30:0] addW_838;
wire [4:0] slice_1027;
wire [14:0] mul4_1216;
wire [14:0] mulnw_1405;
wire [23:0] addW_1594;
wire [19:0] add_1783;
wire [9:0] mulnw_1972;
wire [8:0] mulnw_144;
wire [31:0] addW_333;
wire [22:0] addW_522;
wire [6:0] slice_711;
wire [8:0] mulnw_900;
wire [22:0] concat_1089;
wire [19:0] addW_1278;
wire [9:0] mulnw_1467;
wire [17:0] slice_1656;
wire [13:0] mul_1845;
wire [9:0] slice_206;
wire [9:0] mul_395;
wire [44:0] concat_584;
wire [11:0] addW_773;
wire [21:0] concat_962;
wire [15:0] mul_1151;
wire [63:0] subW_1340;
wire [14:0] concat_1529;
wire [5:0] slice_1718;
wire [28:0] lsl_1907;
wire [23:0] add_79;
wire [9:0] slice_268;
wire [14:0] mulnw_457;
wire [9:0] mul_646;
wire [58:0] concat_835;
wire [4:0] slice_1024;
wire [6:0] slice_1213;
wire [29:0] add_1402;
wire [14:0] mul4_1591;
wire [15:0] lsl_1780;
wire [18:0] lsl_1969;
wire [16:0] add_330;
wire [13:0] mul_519;
wire [6:0] slice_708;
wire [18:0] lsl_897;
wire [6:0] slice_1086;
wire [11:0] mul_1275;
wire [18:0] lsl_1464;
wire [4:0] slice_1653;
wire [14:0] mulnw_1842;
wire [28:0] slice_14;
wire [9:0] slice_203;
wire [9:0] mulnw_392;
wire [6:0] slice_581;
wire [14:0] concat_770;
wire [11:0] addW_959;
wire [28:0] slice_1148;
wire [44:0] addW_1337;
wire [4:0] slice_1526;
wire [87:0] concat_1715;
wire [23:0] add_1904;
wire [15:0] add_76;
wire [4:0] slice_265;
wire [29:0] concat_454;
wire [4:0] slice_643;
wire [42:0] subW_832;
wire [39:0] concat_1021;
wire [6:0] slice_1210;
wire [22:0] lsl_1399;
wire [13:0] mul_1588;
wire [9:0] mulnw_1777;
wire [30:0] concat_1966;
wire [17:0] mul_138;
wire [10:0] add_327;
wire [13:0] mul_516;
wire [14:0] slice_705;
wire [19:0] add_894;
wire [7:0] slice_1083;
wire [11:0] mul_1272;
wire [30:0] concat_1461;
wire [9:0] mul_1650;
wire [14:0] mulnw_1839;
wire [17:0] slice_200;
wire [18:0] lsl_389;
wire [13:0] mul_578;
wire [4:0] slice_767;
wire [14:0] concat_956;
wire [14:0] slice_1145;
wire [40:0] concat_1334;
wire [4:0] slice_1523;
wire [17:0] slice_1712;
wire [15:0] add_1901;
wire [28:0] lsl_73;
wire [55:0] slice_262;
wire [15:0] addW_451;
wire [4:0] slice_640;
wire [8:0] slice_829;
wire [17:0] slice_1018;
wire [14:0] slice_1207;
wire [13:0] mulnw_1396;
wire [15:0] mul_1585;
wire [8:0] mulnw_1774;
wire [8:0] slice_1963;
wire [21:0] concat_135;
wire [4:0] slice_324;
wire [13:0] mul_513;
wire [112:0] slice_702;
wire [15:0] lsl_891;
wire [7:0] slice_1080;
wire [11:0] mul_1269;
wire [8:0] slice_1458;
wire [4:0] slice_1647;
wire [29:0] concat_1836;
wire [17:0] slice_197;
wire [30:0] concat_386;
wire [6:0] slice_575;
wire [4:0] slice_764;
wire [4:0] slice_953;
wire [172:0] concat_1142;
wire [20:0] addW_1331;
wire [4:0] slice_1520;
wire [41:0] subW_1709;
wire [28:0] lsl_1898;
wire [23:0] add_70;
wire [27:0] slice_259;
wire [20:0] concat_448;
wire [9:0] slice_637;
wire [19:0] add_826;
wire [4:0] slice_1015;
wire [14:0] slice_1204;
wire [44:0] concat_1393;
wire [28:0] slice_1582;
wire [16:0] add_1771;
wire [4:0] slice_1960;
wire [11:0] addW_132;
wire [3:0] slice_321;
wire [6:0] slice_510;
wire [28:0] slice_699;
wire [4:0] slice_888;
wire [86:0] concat_1077;
wire [30:0] addW_1266;
wire [4:0] slice_1455;
wire [4:0] slice_1644;
wire [15:0] addW_1833;
wire [19:0] addW_194;
wire [8:0] slice_383;
wire [6:0] slice_572;
wire [4:0] slice_761;
wire [4:0] slice_950;
wire [27:0] slice_1139;
wire [9:0] mul_1328;
wire [43:0] concat_1517;
wire [31:0] addW_1706;
wire [13:0] slice_1895;
wire [15:0] add_67;
wire [63:0] subW_256;
wire [6:0] slice_445;
wire [9:0] slice_634;
wire [15:0] lsl_823;
wire [9:0] mul_1012;
wire [13:0] slice_1201;
wire [6:0] slice_1390;
wire [14:0] slice_1579;
wire [10:0] add_1768;
wire [9:0] mul_1957;
wire [14:0] concat_129;
wire [9:0] mul_318;
wire [6:0] slice_507;
wire [229:0] concat_696;
wire [8:0] mulnw_885;
wire [17:0] slice_1074;
wire [30:0] addW_1263;
wire [9:0] mul_1452;
wire [9:0] slice_1641;
wire [20:0] concat_1830;
wire [11:0] mul_191;
wire [4:0] slice_380;
wire [13:0] slice_569;
wire [59:0] concat_758;
wire [4:0] slice_947;
wire [60:0] subW_1136;
wire [8:0] mulnw_1325;
wire [17:0] slice_1514;
wire [16:0] add_1703;
wire [22:0] addW_1892;
wire [28:0] lsl_64;
wire [44:0] addW_253;
wire [6:0] slice_442;
wire [17:0] slice_631;
wire [9:0] mulnw_820;
wire [4:0] slice_1009;
wire [29:0] add_1198;
wire [13:0] mul_1387;
wire [116:0] concat_1576;
wire [8:0] mulnw_1765;
wire [4:0] slice_1954;
wire [4:0] slice_126;
wire [9:0] mulnw_315;
wire [14:0] mul4_504;
wire [120:0] subW_693;
wire [8:0] slice_882;
wire [41:0] subW_1071;
wire [59:0] concat_1260;
wire [4:0] slice_1449;
wire [9:0] slice_1638;
wire [6:0] slice_1827;
wire [11:0] mul_188;
wire [9:0] mul_377;
wire [30:0] concat_566;
wire [30:0] addW_755;
wire [39:0] concat_944;
wire [45:0] addW_1133;
wire [18:0] lsl_1322;
wire [5:0] slice_1511;
wire [10:0] add_1700;
wire [13:0] mul_1889;
wire [44:0] concat_61;
wire [40:0] concat_250;
wire [13:0] slice_439;
wire [17:0] slice_628;
wire [8:0] mulnw_817;
wire [4:0] slice_1006;
wire [22:0] lsl_1195;
wire [6:0] slice_1384;
wire [64:0] subW_1573;
wire [3:0] slice_1762;
wire [4:0] slice_1951;
wire [4:0] slice_123;
wire [18:0] lsl_312;
wire [6:0] slice_501;
wire [28:0] slice_690;
wire [8:0] slice_879;
wire [31:0] addW_1068;
wire [30:0] addW_1257;
wire [4:0] slice_1446;
wire [13:0] slice_1635;
wire [6:0] slice_1824;
wire [11:0] mul_185;
wire [4:0] slice_374;
wire [16:0] addW_563;
wire [13:0] mul_752;
wire [17:0] slice_941;
wire [23:0] add_1130;
wire [19:0] add_1319;
wire [11:0] mul_1508;
wire [4:0] slice_1697;
wire [13:0] mul_1886;
wire [29:0] concat_58;
wire [20:0] addW_247;
wire [23:0] addW_436;
wire [19:0] addW_625;
wire [16:0] add_814;
wire [9:0] slice_1003;
wire [14:0] mulnw_1192;
wire [6:0] slice_1381;
wire [17:0] slice_1570;
wire [17:0] mul_1759;
wire [9:0] slice_1948;
wire [4:0] slice_120;
wire [30:0] concat_309;
wire [6:0] slice_498;
wire [63:0] subW_687;
wire [16:0] addW_876;
wire [16:0] add_1065;
wire [13:0] mul_1254;
wire [9:0] slice_1443;
wire [29:0] add_1632;
wire [13:0] slice_1821;
wire [343:0] addW_2010;
wire [30:0] addW_182;
wire [4:0] slice_371;
wire [22:0] concat_560;
wire [13:0] mulnw_749;
wire [4:0] slice_938;
wire [15:0] add_1127;
wire [15:0] lsl_1316;
wire [5:0] slice_1505;
wire [3:0] slice_1694;
wire [13:0] mul_1883;
wire [15:0] addW_55;
wire [9:0] mul_244;
wire [14:0] mul4_433;
wire [11:0] mul_622;
wire [10:0] add_811;
wire [9:0] slice_1000;
wire [29:0] add_1189;
wire [13:0] slice_1378;
wire [41:0] subW_1567;
wire [21:0] concat_1756;
wire [9:0] slice_1945;
wire [8:0] slice_306;
wire [14:0] slice_495;
wire [44:0] addW_684;
wire [9:0] mul_873;
wire [10:0] add_1062;
wire [13:0] mulnw_1251;
wire [9:0] slice_1440;
wire [22:0] lsl_1629;
wire [23:0] addW_1818;
wire [231:0] concat_2007;
wire [30:0] addW_179;
wire [9:0] slice_368;
wire [6:0] slice_557;
wire [14:0] mulnw_746;
wire [9:0] mul_935;
wire [28:0] lsl_1124;
wire [4:0] slice_1313;
wire [5:0] slice_1502;
wire [9:0] mul_1691;
wire [6:0] slice_1880;
wire [8:0] mulnw_241;
wire [13:0] mul_430;
wire [11:0] mul_619;
wire [8:0] mulnw_808;
wire [17:0] slice_997;
wire [22:0] lsl_1186;
wire [30:0] concat_1375;
wire [31:0] addW_1564;
wire [11:0] addW_1753;
wire [17:0] slice_1942;
wire [17:0] slice_114;
wire [4:0] slice_303;
wire [7:0] slice_492;
wire [40:0] concat_681;
wire [9:0] mul_870;
wire [4:0] slice_1059;
wire [14:0] mulnw_1248;
wire [17:0] slice_1437;
wire [14:0] mulnw_1626;
wire [14:0] mul4_1815;
wire [120:0] subW_2004;
wire [87:0] concat_176;
wire [9:0] slice_365;
wire [7:0] slice_554;
wire [13:0] mul_743;
wire [4:0] slice_932;
wire [23:0] add_1121;
wire [8:0] mulnw_1310;
wire [11:0] slice_1499;
wire [9:0] mulnw_1688;
wire [6:0] slice_1877;
wire [13:0] mul_49;
wire [18:0] lsl_238;
wire [15:0] mul_427;
wire [11:0] mul_616;
wire [3:0] slice_805;
wire [41:0] subW_994;
wire [13:0] mulnw_1183;
wire [16:0] addW_1372;
wire [16:0] add_1561;
wire [14:0] concat_1750;
wire [17:0] slice_1939;
wire [17:0] slice_111;
wire [9:0] mul_300;
wire [58:0] addW_489;
wire [20:0] addW_678;
wire [9:0] mul_867;
wire [3:0] slice_1056;
wire [13:0] mul_1245;
wire [17:0] slice_1434;
wire [29:0] add_1623;
wire [13:0] mul_1812;
wire [28:0] slice_2001;
wire [58:0] concat_173;
wire [17:0] slice_362;
wire [7:0] slice_551;
wire [14:0] mulnw_740;
wire [4:0] slice_929;
wire [15:0] add_1118;
wire [8:0] slice_1307;
wire [11:0] slice_1496;
wire [18:0] lsl_1685;
wire [14:0] mul4_1874;
wire [13:0] mul_46;
wire [19:0] add_235;
wire [29:0] addW_424;
wire [30:0] addW_613;
wire [17:0] mul_802;
wire [31:0] addW_991;
wire [44:0] concat_1180;
wire [22:0] concat_1369;
wire [10:0] add_1558;
wire [4:0] slice_1747;
wire [19:0] addW_1936;
wire [21:0] concat_108;
wire [4:0] slice_297;
wire [172:0] concat_486;
wire [9:0] mul_675;
wire [19:0] addW_864;
wire [9:0] mul_1053;
wire [14:0] mulnw_1242;
wire [16:0] addW_1431;
wire [22:0] lsl_1620;
wire [15:0] mul_1809;
wire [63:0] subW_1998;
wire [42:0] subW_170;
wire [17:0] slice_359;
wire [59:0] concat_548;
wire [14:0] mulnw_737;
wire [9:0] slice_926;
wire [28:0] lsl_1115;
wire [8:0] slice_1304;
wire [27:0] slice_1493;
wire [30:0] concat_1682;
wire [6:0] slice_1871;
wire [6:0] slice_43;
wire [15:0] lsl_232;
wire [29:0] addW_421;
wire [30:0] addW_610;
wire [21:0] concat_799;
wire [16:0] add_988;
wire [6:0] slice_1177;
wire [6:0] slice_1366;
wire [4:0] slice_1555;
wire [4:0] slice_1744;
wire [11:0] mul_1933;
wire [11:0] addW_105;
wire [4:0] slice_294;
wire [115:0] concat_483;
wire [8:0] mulnw_672;
wire [19:0] addW_861;
wire [9:0] mulnw_1050;
wire [14:0] mulnw_1239;
wire [9:0] mul_1428;
wire [13:0] mulnw_1617;
wire [28:0] slice_1806;
wire [44:0] addW_1995;
wire [8:0] slice_167;
wire [16:0] addW_356;
wire [30:0] addW_545;
wire [29:0] concat_734;
wire [4:0] slice_923;
wire [13:0] slice_1112;
wire [16:0] addW_1301;
wire [40:0] addW_1490;
wire [8:0] slice_1679;
wire [6:0] slice_1868;
wire [30:0] concat_40;
wire [4:0] slice_229;
wire [27:0] slice_418;
wire [28:0] slice_607;
wire [11:0] addW_796;
wire [10:0] add_985;
wire [13:0] mul_1174;
wire [7:0] slice_1363;
wire [3:0] slice_1552;
wire [4:0] slice_1741;
wire [11:0] mul_1930;
wire [9:0] slice_291;
wire [61:0] subW_480;
wire [18:0] lsl_669;
wire [35:0] mul_858;
wire [18:0] lsl_1047;
wire [29:0] concat_1236;
wire [9:0] mul_1425;
wire [44:0] concat_1614;
wire [14:0] slice_1803;
wire [40:0] concat_1992;
wire [19:0] add_164;
wire [9:0] mul_353;
wire [13:0] mul_542;
wire [15:0] addW_731;
wire [55:0] slice_920;
wire [22:0] addW_1109;
wire [9:0] mul_1298;
wire [40:0] concat_1487;
wire [4:0] slice_1676;
wire [14:0] slice_1865;
wire [16:0] addW_37;
wire [8:0] mulnw_226;
wire [40:0] addW_415;
wire [45:0] addW_604;
wire [14:0] concat_793;
wire [4:0] slice_982;
wire [6:0] slice_1171;
wire [56:0] slice_1360;
wire [9:0] mul_1549;
wire [43:0] concat_1738;
wire [11:0] mul_1927;
wire [9:0] mul_99;
wire [9:0] slice_288;
wire [13:0] slice_477;
wire [19:0] add_666;
wire [25:0] concat_855;
wire [30:0] concat_1044;
wire [15:0] addW_1233;
wire [9:0] mul_1422;
wire [6:0] slice_1611;
wire [20:0] addW_1989;
wire [15:0] lsl_161;
wire [9:0] mul_350;
wire [13:0] mulnw_539;
wire [20:0] concat_728;
wire [88:0] addW_917;
wire [13:0] mul_1106;
wire [9:0] mul_1295;
wire [20:0] addW_1484;
wire [9:0] mul_1673;
wire [14:0] slice_1862;
wire [8:0] slice_223;
wire [40:0] concat_412;
wire [23:0] add_601;
wire [4:0] slice_790;
wire [3:0] slice_979;
wire [6:0] slice_1168;
wire [14:0] slice_1357;
wire [9:0] mulnw_1546;
wire [17:0] slice_1735;
wire [30:0] addW_1924;
wire [17:0] slice_285;
wire [29:0] add_474;
wire [15:0] lsl_663;
wire [13:0] addW_852;
wire [8:0] slice_1041;
wire [20:0] concat_1230;
wire [27:0] slice_1419;
wire [13:0] mul_1608;
wire [116:0] concat_1797;
wire [9:0] mul_1986;
wire [9:0] mulnw_158;
wire [9:0] mul_347;
wire [14:0] mulnw_536;
wire [6:0] slice_725;
wire [62:0] concat_914;
wire [13:0] mul_1103;
wire [9:0] mul_1292;
wire [9:0] mul_1481;
wire [4:0] slice_1670;
wire [13:0] slice_1859;
wire [8:0] slice_220;
wire [20:0] addW_409;
wire [15:0] add_598;
wire [4:0] slice_787;
wire [9:0] mul_976;
wire [13:0] slice_1165;
wire [114:0] addW_1354;
wire [18:0] lsl_1543;
wire [5:0] slice_1732;
wire [30:0] addW_1921;
wire [9:0] slice_93;
wire [17:0] slice_282;
wire [22:0] lsl_471;
wire [4:0] slice_660;
wire [17:0] concat_849;
wire [4:0] slice_1038;
wire [6:0] slice_1227;
wire [27:0] slice_1416;
wire [6:0] slice_1605;
wire [64:0] subW_1794;
wire [8:0] mulnw_1983;
wire [8:0] mulnw_155;
wire [27:0] slice_344;
wire [13:0] mul_533;
wire [6:0] slice_722;
wire [42:0] subW_911;
wire [13:0] mul_1100;
wire [19:0] addW_1289;
wire [8:0] mulnw_1478;
wire [4:0] slice_1667;
wire [29:0] add_1856;
wire [6:0] slice_28;
wire [16:0] addW_217;
wire [9:0] mul_406;
wire [28:0] lsl_595;
wire [4:0] slice_784;
wire [9:0] mulnw_973;
wire [30:0] concat_1162;
wire [342:0] concat_1351;
wire [30:0] concat_1540;
wire [11:0] mul_1729;
wire [59:0] concat_1918;
wire [16:0] addW_279;
wire [14:0] mulnw_468;
wire [8:0] mulnw_657;
wire [5:0] slice_846;
wire [9:0] mul_1035;
wire [6:0] slice_1224;
wire [45:0] addW_1413;
wire [6:0] slice_1602;
wire [17:0] slice_1791;
wire [18:0] lsl_1980;
wire [16:0] add_152;
wire [27:0] slice_341;
wire [14:0] mulnw_530;
wire [13:0] slice_719;
wire [8:0] slice_908;
wire [6:0] slice_1097;
wire [19:0] addW_1286;
wire [18:0] lsl_1475;
wire [9:0] slice_1664;
wire [22:0] lsl_1853;
wire [15:0] mul_25;
wire [9:0] mul_214;
wire [8:0] mulnw_403;
wire [23:0] add_592;
wire [39:0] concat_781;
wire [18:0] lsl_970;
wire [16:0] addW_1159;
wire [55:0] slice_1348;
wire [8:0] slice_1537;
wire [5:0] slice_1726;
wire [30:0] addW_1915;
wire [27:0] slice_87;
wire [9:0] mul_276;
wire [29:0] add_465;
wire [8:0] slice_654;
wire [5:0] slice_843;
wire [4:0] slice_1032;
wire [13:0] slice_1221;
wire [23:0] add_1410;
wire [13:0] slice_1599;
wire [41:0] subW_1788;
wire [19:0] add_1977;
wire [10:0] add_149;
wire [40:0] addW_338;
wire [14:0] mulnw_527;
wire [23:0] addW_716;
wire [19:0] add_905;
wire [6:0] slice_1094;
wire [35:0] mul_1283;
wire [19:0] add_1472;
wire [9:0] slice_1661;
wire [14:0] mulnw_1850;
wire [28:0] slice_22;
wire [9:0] mul_211;
wire [18:0] lsl_400;
wire [15:0] add_589;
wire [17:0] slice_778;
wire [30:0] concat_967;
wire [22:0] concat_1156;
wire [119:0] subW_1345;
wire [4:0] slice_1534;
wire [5:0] slice_1723;
wire [13:0] mul_1912;
wire [59:0] concat_84;
wire [9:0] mul_273;
wire [22:0] lsl_462;
wire [8:0] slice_651;
wire [5:0] slice_840;
wire [4:0] slice_1029;
wire [23:0] addW_1218;
wire [15:0] add_1407;
wire [30:0] concat_1596;
wire [31:0] addW_1785;
wire [15:0] lsl_1974;
wire [8:0] mulnw_146;
wire [40:0] concat_335;
wire [29:0] concat_524;
wire [14:0] mul4_713;
wire [15:0] lsl_902;
wire [14:0] mul4_1091;
wire [25:0] concat_1280;
wire [15:0] lsl_1469;
wire [17:0] slice_1658;
wire [29:0] add_1847;
wire [9:0] mul_208;
wire [19:0] add_397;
wire [28:0] lsl_586;
wire [4:0] slice_775;
wire [8:0] slice_964;
wire [6:0] slice_1153;
wire [89:0] addW_1342;
wire [9:0] mul_1531;
wire [11:0] slice_1720;
wire [13:0] mulnw_1909;
wire [30:0] addW_81;
wire [9:0] mul_270;
wire [13:0] mulnw_459;
wire [16:0] addW_648;
wire [87:0] concat_837;
wire [9:0] slice_1026;
wire [14:0] mul4_1215;
wire [28:0] lsl_1404;
wire [16:0] addW_1593;
wire [16:0] add_1782;
wire [4:0] slice_1971;
wire [3:0] slice_143;
wire [20:0] addW_332;
wire [15:0] addW_521;
wire [13:0] mul_710;
wire [9:0] mulnw_899;
wire [6:0] slice_1088;
wire [13:0] addW_1277;
wire [4:0] slice_1466;
wire [17:0] slice_1655;
wire [22:0] lsl_1844;
wire [14:0] slice_16;
wire [19:0] addW_205;
wire [15:0] lsl_394;
wire [13:0] slice_583;
wire [9:0] mul_772;
wire [4:0] slice_961;
wire [7:0] slice_1150;
wire [62:0] concat_1339;
wire [4:0] slice_1528;
wire [11:0] slice_1717;
wire [14:0] mulnw_1906;
wire [13:0] mul_78;
wire [27:0] slice_267;
wire [44:0] concat_456;
wire [9:0] mul_645;
wire [17:0] slice_834;
wire [9:0] slice_1023;
wire [13:0] mul_1212;
wire [23:0] add_1401;
wire [22:0] concat_1590;
wire [10:0] add_1779;
wire [8:0] mulnw_1968;
wire [30:0] concat_140;
wire [9:0] mul_329;
wire [20:0] concat_518;
wire [15:0] mul_707;
wire [8:0] mulnw_896;
wire [6:0] slice_1085;
wire [17:0] concat_1274;
wire [8:0] mulnw_1463;
wire [16:0] addW_1652;
wire [13:0] mulnw_1841;
wire [19:0] addW_202;
wire [4:0] slice_391;
wire [22:0] addW_580;
wire [4:0] slice_769;
wire [9:0] mul_958;
wire [58:0] addW_1147;
wire [42:0] subW_1336;
wire [4:0] slice_1525;
wire [27:0] slice_1714;
wire [13:0] mul_1903;
wire [13:0] mulnw_75;
wire [9:0] slice_264;
wire [6:0] slice_453;
wire [9:0] mul_642;
wire [41:0] subW_831;
wire [17:0] slice_1020;
wire [15:0] mul_1209;
wire [15:0] add_1398;
wire [6:0] slice_1587;
wire [4:0] slice_1776;
wire [8:0] slice_1965;
wire [8:0] slice_137;
wire [8:0] mulnw_326;
wire [6:0] slice_515;
wire [28:0] slice_704;
wire [16:0] add_893;
wire [14:0] slice_1082;
wire [5:0] slice_1271;
wire [8:0] slice_1460;
wire [9:0] mul_1649;
wire [44:0] concat_1838;
wire [35:0] mul_199;
wire [8:0] mulnw_388;
wire [13:0] mul_577;
wire [4:0] slice_766;
wire [4:0] slice_955;
wire [28:0] slice_1144;
wire [8:0] slice_1333;
wire [9:0] slice_1522;
wire [40:0] addW_1711;
wire [14:0] mulnw_1900;
wire [14:0] mulnw_72;
wire [13:0] mul_450;
wire [9:0] mul_639;
wire [31:0] addW_828;
wire [17:0] slice_1017;
wire [28:0] slice_1206;
wire [28:0] lsl_1395;
wire [7:0] slice_1584;
wire [3:0] slice_1773;
wire [8:0] slice_1962;
wire [4:0] slice_134;
wire [18:0] lsl_323;
wire [6:0] slice_512;
wire [7:0] slice_701;
wire [10:0] add_890;
wire [14:0] slice_1079;
wire [5:0] slice_1268;
wire [8:0] slice_1457;
wire [9:0] mul_1646;
wire [6:0] slice_1835;
wire [25:0] concat_196;
wire [8:0] slice_385;
wire [13:0] mul_574;
wire [9:0] slice_763;
wire [4:0] slice_952;
wire [55:0] slice_1141;
wire [19:0] add_1330;
wire [9:0] slice_1519;
wire [40:0] concat_1708;
wire [14:0] mulnw_1897;
wire [13:0] mul_69;
wire [88:0] addW_258;
wire [6:0] slice_447;
wire [19:0] addW_636;
wire [16:0] add_825;
wire [16:0] addW_1014;
wire [28:0] slice_1203;
wire [13:0] slice_1392;
wire [56:0] slice_1581;
wire [9:0] mul_1770;
wire [16:0] addW_1959;
wire [9:0] mul_131;
wire [19:0] add_320;
wire [13:0] slice_509;
wire [56:0] slice_698;
wire [8:0] mulnw_887;
wire [27:0] slice_1076;
wire [5:0] slice_1265;
wire [16:0] addW_1454;
wire [9:0] mul_1643;
wire [13:0] mul_1832;
wire [13:0] addW_193;
wire [8:0] slice_382;
wire [13:0] mul_571;
wire [9:0] slice_760;
wire [9:0] slice_949;
wire [87:0] addW_1138;
wire [15:0] lsl_1327;
wire [17:0] slice_1516;
wire [20:0] addW_1705;
wire [29:0] concat_1894;
wire [14:0] mulnw_66;
wire [62:0] concat_255;
wire [6:0] slice_444;
wire [19:0] addW_633;
wire [10:0] add_822;
wire [9:0] mul_1011;
wire [45:0] addW_1200;
wire [22:0] addW_1389;
wire [28:0] slice_1578;
wire [9:0] mulnw_1767;
wire [9:0] mul_1956;
wire [4:0] slice_128;
wire [15:0] lsl_317;
wire [23:0] addW_506;
wire [55:0] slice_695;
wire [3:0] slice_884;
wire [40:0] addW_1073;
wire [88:0] concat_1262;
wire [9:0] mul_1451;
wire [27:0] slice_1640;
wire [6:0] slice_1829;
wire [17:0] concat_190;
wire [16:0] addW_379;
wire [6:0] slice_568;
wire [13:0] slice_757;
wire [9:0] slice_946;
wire [59:0] concat_1135;
wire [9:0] mulnw_1324;
wire [17:0] slice_1513;
wire [9:0] mul_1702;
wire [15:0] addW_1891;
wire [14:0] mulnw_63;
wire [42:0] subW_252;
wire [13:0] slice_441;
wire [35:0] mul_630;
wire [4:0] slice_819;
wire [9:0] mul_1008;
wire [23:0] add_1197;
wire [13:0] mul_1386;
wire [27:0] slice_1575;
wire [18:0] lsl_1764;
wire [9:0] mul_1953;
wire [4:0] slice_125;
wire [4:0] slice_314;
wire [14:0] mul4_503;
wire [119:0] subW_692;
wire [17:0] mul_881;
wire [40:0] concat_1070;
wire [13:0] slice_1259;
wire [9:0] mul_1448;
wire [27:0] slice_1637;
wire [6:0] slice_1826;
wire [5:0] slice_187;
wire [9:0] mul_376;
wire [6:0] slice_565;
wire [29:0] add_754;
wire [17:0] slice_943;
wire [30:0] addW_1132;
wire [8:0] mulnw_1321;
wire [19:0] addW_1510;
wire [8:0] mulnw_1699;
wire [20:0] concat_1888;
wire [13:0] slice_60;
wire [8:0] slice_249;
wire [30:0] concat_438;
wire [25:0] concat_627;
wire [3:0] slice_816;
wire [9:0] mul_1005;
wire [15:0] add_1194;
wire [13:0] mul_1383;
wire [63:0] subW_1572;
wire [30:0] concat_1761;
wire [9:0] mul_1950;
wire [9:0] slice_122;
wire [8:0] mulnw_311;
wire [13:0] mul_500;
wire [89:0] addW_689;
wire [21:0] concat_878;
wire [20:0] addW_1067;
wire [29:0] add_1256;
wire [9:0] mul_1445;
wire [45:0] addW_1634;
wire [13:0] slice_1823;
wire [456:0] concat_2012;
wire [5:0] slice_184;
wire [9:0] mul_373;
wire [14:0] mul4_562;
wire [22:0] lsl_751;
wire [17:0] slice_940;
wire [13:0] mul_1129;
wire [16:0] add_1318;
wire [11:0] mul_1507;
wire [18:0] lsl_1696;
wire [6:0] slice_1885;
wire [6:0] slice_57;
wire [19:0] add_246;
wire [16:0] addW_435;
wire [13:0] addW_624;
wire [9:0] mul_813;
wire [27:0] slice_1002;
wire [28:0] lsl_1191;
wire [13:0] mul_1380;
wire [44:0] addW_1569;
wire [8:0] slice_1758;
wire [19:0] addW_1947;
wire [9:0] slice_119;
wire [8:0] slice_308;
wire [15:0] mul_497;
wire [62:0] concat_686;
wire [11:0] addW_875;
wire [9:0] mul_1064;
wire [22:0] lsl_1253;
wire [19:0] addW_1442;
wire [23:0] add_1631;
wire [30:0] concat_1820;
wire [233:0] subW_2009;
wire [5:0] slice_181;
wire [9:0] mul_370;
wire [6:0] slice_559;
wire [14:0] mulnw_748;
wire [16:0] addW_937;
wire [13:0] mulnw_1126;
wire [10:0] add_1315;
wire [11:0] mul_1504;
wire [19:0] add_1693;
wire [6:0] slice_1882;
wire [13:0] mul_54;
wire [15:0] lsl_243;
wire [22:0] concat_432;
wire [17:0] concat_621;
wire [9:0] mulnw_810;
wire [27:0] slice_999;
wire [23:0] add_1188;
wire [6:0] slice_1377;
wire [40:0] concat_1566;
wire [4:0] slice_1755;
wire [19:0] addW_1944;
wire [8:0] slice_305;
wire [28:0] slice_494;
wire [42:0] subW_683;
wire [14:0] concat_872;
wire [8:0] mulnw_1061;
wire [14:0] mulnw_1250;
wire [19:0] addW_1439;
wire [15:0] add_1628;
wire [16:0] addW_1817;
wire [56:0] slice_2006;
wire [19:0] addW_367;
wire [6:0] slice_556;
wire [29:0] add_745;
wire [9:0] mul_934;
wire [14:0] mulnw_1123;
wire [8:0] mulnw_1312;
wire [11:0] mul_1501;
wire [15:0] lsl_1690;
wire [13:0] slice_1879;
wire [20:0] concat_51;
wire [9:0] mulnw_240;
wire [6:0] slice_429;
wire [5:0] slice_618;
wire [18:0] lsl_807;
wire [40:0] addW_996;
wire [15:0] add_1185;
wire [6:0] slice_1374;
wire [20:0] addW_1563;
wire [9:0] mul_1752;
wire [35:0] mul_1941;
wire [16:0] addW_302;
wire [14:0] slice_491;
wire [8:0] slice_680;
wire [4:0] slice_869;
wire [18:0] lsl_1058;
wire [29:0] add_1247;
wire [35:0] mul_1436;
wire [28:0] lsl_1625;
wire [22:0] concat_1814;
wire [119:0] subW_2003;
wire [27:0] slice_175;
wire [19:0] addW_364;
wire [14:0] slice_553;
wire [22:0] lsl_742;
wire [9:0] mul_931;
wire [13:0] mul_1120;
wire [3:0] slice_1309;
wire [30:0] addW_1498;
wire [4:0] slice_1687;
wire [23:0] addW_1876;
wire [6:0] slice_48;
wire [8:0] mulnw_237;
wire [7:0] slice_426;
wire [5:0] slice_615;
wire [30:0] concat_804;
wire [40:0] concat_993;
wire [28:0] lsl_1182;
wire [14:0] mul4_1371;
wire [9:0] mul_1560;
wire [4:0] slice_1749;
wire [25:0] concat_1938;
wire [17:0] slice_110;
wire [9:0] mul_299;
wire [19:0] add_677;
wire [4:0] slice_866;
wire [19:0] add_1055;
wire [22:0] lsl_1244;
wire [21:0] concat_1433;
wire [23:0] add_1622;
wire [6:0] slice_1811;
wire [89:0] addW_2000;
wire [17:0] slice_172;
wire [35:0] mul_361;
wire [14:0] slice_550;
wire [13:0] mulnw_739;
wire [9:0] mul_928;
wire [14:0] mulnw_1117;
wire [17:0] mul_1306;
wire [30:0] addW_1495;
wire [8:0] mulnw_1684;
wire [14:0] mul4_1873;
wire [6:0] slice_45;
wire [16:0] add_234;
wire [7:0] slice_423;
wire [5:0] slice_612;
wire [8:0] slice_801;
wire [20:0] addW_990;
wire [13:0] slice_1179;
wire [6:0] slice_1368;
wire [8:0] mulnw_1557;
wire [4:0] slice_1746;
wire [13:0] addW_1935;
wire [4:0] slice_107;
wire [9:0] mul_296;
wire [55:0] slice_485;
wire [15:0] lsl_674;
wire [4:0] slice_863;
wire [15:0] lsl_1052;
wire [13:0] mulnw_1241;
wire [11:0] addW_1430;
wire [15:0] add_1619;
wire [7:0] slice_1808;
wire [62:0] concat_1997;
wire [41:0] subW_169;
wire [21:0] concat_358;
wire [13:0] slice_547;
wire [44:0] concat_736;
wire [27:0] slice_925;
wire [14:0] mulnw_1114;
wire [21:0] concat_1303;
wire [58:0] concat_1492;
wire [8:0] slice_1681;
wire [13:0] mul_1870;
wire [13:0] slice_42;
wire [10:0] add_231;
wire [4:0] slice_798;
wire [9:0] mul_987;
wire [22:0] addW_1176;
wire [6:0] slice_1365;
wire [18:0] lsl_1554;
wire [9:0] slice_1743;
wire [17:0] concat_1932;
wire [9:0] mul_104;
wire [9:0] mul_293;
wire [27:0] slice_482;
wire [9:0] mulnw_671;
wire [43:0] concat_860;
wire [4:0] slice_1049;
wire [44:0] concat_1238;
wire [14:0] concat_1427;
wire [28:0] lsl_1616;
wire [58:0] addW_1805;
wire [42:0] subW_1994;
wire [31:0] addW_166;
wire [11:0] addW_355;
wire [29:0] add_544;
wire [6:0] slice_733;
wire [9:0] slice_922;
wire [29:0] concat_1111;
wire [11:0] addW_1300;
wire [42:0] subW_1489;
wire [8:0] slice_1678;
wire [15:0] mul_1867;
wire [6:0] slice_39;
wire [8:0] mulnw_228;
wire [58:0] concat_417;
wire [59:0] concat_606;
wire [9:0] mul_795;
wire [8:0] mulnw_984;
wire [13:0] mul_1173;
wire [14:0] slice_1362;
wire [19:0] add_1551;
wire [9:0] slice_1740;
wire [5:0] slice_1929;
wire [14:0] concat_101;
wire [19:0] addW_290;
wire [60:0] subW_479;
wire [8:0] mulnw_668;
wire [17:0] slice_857;
wire [8:0] mulnw_1046;
wire [6:0] slice_1235;
wire [4:0] slice_1424;
wire [13:0] slice_1613;
wire [28:0] slice_1802;
wire [8:0] slice_1991;
wire [16:0] add_163;
wire [14:0] concat_352;
wire [22:0] lsl_541;
wire [13:0] mul_730;
wire [116:0] concat_919;
wire [15:0] addW_1108;
wire [14:0] concat_1297;
wire [8:0] slice_1486;
wire [16:0] addW_1675;
wire [28:0] slice_1864;
wire [14:0] mul4_36;
wire [3:0] slice_225;
wire [42:0] subW_414;
wire [30:0] addW_603;
wire [4:0] slice_792;
wire [18:0] lsl_981;
wire [13:0] mul_1170;
wire [114:0] addW_1359;
wire [15:0] lsl_1548;
wire [17:0] slice_1737;
wire [5:0] slice_1926;
wire [4:0] slice_98;
wire [19:0] addW_287;
wire [45:0] addW_476;
wire [16:0] add_665;
wire [5:0] slice_854;
wire [8:0] slice_1043;
wire [13:0] mul_1232;
wire [4:0] slice_1421;
wire [22:0] addW_1610;
wire [173:0] concat_1799;
wire [19:0] add_1988;
wire [10:0] add_160;
wire [4:0] slice_349;
wire [14:0] mulnw_538;
wire [6:0] slice_727;
wire [64:0] subW_916;
wire [20:0] concat_1105;
wire [4:0] slice_1294;
wire [19:0] add_1483;
wire [9:0] mul_1672;
wire [28:0] slice_1861;
wire [22:0] concat_33;
wire [17:0] mul_222;
wire [8:0] slice_411;
wire [13:0] mul_600;
wire [4:0] slice_789;
wire [19:0] add_978;
wire [13:0] mul_1167;
wire [28:0] slice_1356;
wire [4:0] slice_1545;
wire [17:0] slice_1734;
wire [5:0] slice_1923;
wire [9:0] mul_95;
wire [35:0] mul_284;
wire [23:0] add_473;
wire [10:0] add_662;
wire [11:0] mul_851;
wire [8:0] slice_1040;
wire [6:0] slice_1229;
wire [4:0] slice_1418;
wire [13:0] mul_1607;
wire [27:0] slice_1796;
wire [15:0] lsl_1985;
wire [4:0] slice_157;
wire [4:0] slice_346;
wire [29:0] add_535;
wire [6:0] slice_724;
wire [17:0] slice_913;
wire [6:0] slice_1102;
wire [4:0] slice_1291;
wire [15:0] lsl_1480;
wire [9:0] mul_1669;
wire [45:0] addW_1858;
wire [13:0] mul_30;
wire [21:0] concat_219;
wire [19:0] add_408;
wire [13:0] mulnw_597;
wire [9:0] slice_786;
wire [15:0] lsl_975;
wire [6:0] slice_1164;
wire [8:0] mulnw_1542;
wire [19:0] addW_1731;
wire [88:0] concat_1920;
wire [27:0] slice_92;
wire [21:0] concat_281;
wire [15:0] add_470;
wire [8:0] mulnw_659;
wire [5:0] slice_848;
wire [16:0] addW_1037;
wire [6:0] slice_1226;
wire [59:0] concat_1415;
wire [13:0] mul_1604;
wire [63:0] subW_1793;
wire [9:0] mulnw_1982;
wire [3:0] slice_154;
wire [4:0] slice_343;
wire [22:0] lsl_532;
wire [13:0] slice_721;
wire [41:0] subW_910;
wire [6:0] slice_1099;
wire [4:0] slice_1288;
wire [9:0] mulnw_1477;
wire [9:0] mul_1666;
wire [23:0] add_1855;
wire [11:0] addW_216;
wire [15:0] lsl_405;
wire [14:0] mulnw_594;
wire [9:0] slice_783;
wire [4:0] slice_972;
wire [6:0] slice_1161;
wire [112:0] slice_1350;
wire [8:0] slice_1539;
wire [11:0] mul_1728;
wire [13:0] slice_1917;
wire [9:0] slice_89;
wire [11:0] addW_278;
wire [28:0] lsl_467;
wire [3:0] slice_656;
wire [5:0] slice_845;
wire [9:0] mul_1034;
wire [13:0] slice_1223;
wire [30:0] addW_1412;
wire [13:0] mul_1601;
wire [44:0] addW_1790;
wire [8:0] mulnw_1979;
wire [9:0] mul_151;
wire [58:0] concat_340;
wire [13:0] mulnw_529;
wire [30:0] concat_718;
wire [31:0] addW_907;
wire [13:0] slice_1096;
wire [43:0] concat_1285;
wire [8:0] mulnw_1474;
wire [19:0] addW_1663;
wire [15:0] add_1852;
wire [7:0] slice_24;
wire [14:0] concat_213;
wire [9:0] mulnw_402;
wire [13:0] mul_591;
wire [17:0] slice_780;
wire [8:0] mulnw_969;
wire [14:0] mul4_1158;
wire [173:0] addW_1347;
wire [8:0] slice_1536;
wire [11:0] mul_1725;
wire [29:0] add_1914;
wire [14:0] concat_275;
wire [23:0] add_464;
wire [17:0] mul_653;
wire [11:0] slice_842;
wire [9:0] mul_1031;
wire [30:0] concat_1220;
wire [13:0] mul_1409;
wire [6:0] slice_1598;
wire [40:0] concat_1787;
wire [16:0] add_1976;
wire [9:0] mulnw_148;
wire [42:0] subW_337;
wire [44:0] concat_526;
wire [16:0] addW_715;
wire [16:0] add_904;
wire [23:0] addW_1093;
wire [17:0] slice_1282;
wire [16:0] add_1471;
wire [19:0] addW_1660;
wire [28:0] lsl_1849;
wire [56:0] slice_21;
wire [4:0] slice_210;
wire [8:0] mulnw_399;
wire [14:0] mulnw_588;
wire [17:0] slice_777;
wire [8:0] slice_966;
wire [6:0] slice_1155;
wire [118:0] concat_1344;
wire [16:0] addW_1533;
wire [11:0] mul_1722;
wire [22:0] lsl_1911;
wire [13:0] slice_83;
wire [4:0] slice_272;
wire [15:0] add_461;
wire [21:0] concat_650;
wire [11:0] slice_839;
wire [9:0] mul_1028;
wire [16:0] addW_1217;
wire [13:0] mulnw_1406;
wire [6:0] slice_1595;
wire [20:0] addW_1784;
wire [10:0] add_1973;
wire [18:0] lsl_145;
wire [8:0] slice_334;
wire [6:0] slice_523;
wire [22:0] concat_712;
wire [10:0] add_901;
wire [14:0] mul4_1090;
wire [5:0] slice_1279;
wire [10:0] add_1468;
wire [35:0] mul_1657;
wire [23:0] add_1846;
wire [7:0] slice_18;
wire [4:0] slice_207;
wire [16:0] add_396;
wire [14:0] mulnw_585;
wire [16:0] addW_774;
wire [8:0] slice_963;
wire [6:0] slice_1152;
wire [64:0] subW_1341;
wire [9:0] mul_1530;
wire [30:0] addW_1719;
wire [14:0] mulnw_1908;
wire [29:0] add_80;
wire [4:0] slice_269;
wire [28:0] lsl_458;
wire [11:0] addW_647;
wire [27:0] slice_836;
wire [19:0] addW_1025;
wire [22:0] concat_1214;
wire [14:0] mulnw_1403;
wire [14:0] mul4_1592;
wire [9:0] mul_1781;
wire [8:0] mulnw_1970;
wire [19:0] add_331;
wire [13:0] mul_520;
wire [6:0] slice_709;
wire [4:0] slice_898;
wire [13:0] mul_1087;
wire [11:0] mul_1276;
wire [8:0] mulnw_1465;
wire [21:0] concat_1654;
wire [15:0] add_1843;
wire [4:0] slice_204;
wire [10:0] add_393;
wire [29:0] concat_582;
wire [9:0] mul_771;
wire [16:0] addW_960;
wire [14:0] slice_1149;
wire [17:0] slice_1338;
wire [9:0] mul_1527;
wire [30:0] addW_1716;
wire [29:0] add_1905;
wire [22:0] lsl_77;
wire [55:0] slice_266;
wire [13:0] slice_455;
wire [14:0] concat_644;
wire [40:0] addW_833;
wire [19:0] addW_1022;
wire [6:0] slice_1211;
wire [13:0] mul_1400;
wire [6:0] slice_1589;
wire [8:0] mulnw_1778;
wire [3:0] slice_1967;
wire [8:0] slice_139;
wire [15:0] lsl_328;
wire [6:0] slice_517;
wire [7:0] slice_706;
wire [3:0] slice_895;
wire [15:0] mul_1084;
wire [5:0] slice_1273;
wire [3:0] slice_1462;
wire [11:0] addW_1651;
wire [28:0] lsl_1840;
wire [56:0] slice_12;
wire [43:0] concat_201;
wire [8:0] mulnw_390;
wire [15:0] addW_579;
wire [9:0] mul_768;
wire [9:0] mul_957;
wire [7:0] slice_1146;
wire [41:0] subW_1335;
wire [9:0] mul_1524;
wire [58:0] concat_1713;
wire [22:0] lsl_1902;
wire [14:0] mulnw_74;
wire [27:0] slice_263;
wire [22:0] addW_452;
wire [4:0] slice_641;
wire [40:0] concat_830;
wire [35:0] mul_1019;
wire [7:0] slice_1208;
wire [14:0] mulnw_1397;
wire [6:0] slice_1586;
wire [18:0] lsl_1775;
wire [17:0] mul_1964;
wire [8:0] slice_136;
wire [9:0] mulnw_325;
wire [6:0] slice_514;
wire [56:0] slice_703;
wire [9:0] mul_892;
wire [29:0] addW_1081;
wire [5:0] slice_1270;
wire [17:0] mul_1459;
wire [14:0] concat_1648;
wire [13:0] slice_1837;
wire [112:0] slice_9;
wire [17:0] slice_198;
wire [3:0] slice_387;
wire [20:0] concat_576;
wire [9:0] mul_765;
wire [9:0] mul_954;
wire [58:0] addW_1143;
wire [31:0] addW_1332;
wire [19:0] addW_1521;
wire [42:0] subW_1710;
wire [13:0] mulnw_1899;
wire [29:0] add_71;
wire [116:0] concat_260;
wire [13:0] mul_449;
wire [4:0] slice_638;
wire [20:0] addW_827;
wire [21:0] concat_1016;
wire [7:0] slice_1205;
wire [14:0] mulnw_1394;
wire [14:0] slice_1583;
wire [19:0] add_1772;
wire [21:0] concat_1961;
wire [16:0] addW_133;
wire [8:0] mulnw_322;
wire [13:0] slice_511;
wire [14:0] slice_700;
wire [9:0] mulnw_889;
wire [29:0] addW_1078;
wire [11:0] slice_1267;
wire [21:0] concat_1456;
wire [4:0] slice_1645;
wire [22:0] addW_1834;
wire [5:0] slice_195;
wire [17:0] mul_384;
wire [6:0] slice_573;
wire [27:0] slice_762;
wire [9:0] mul_951;
wire [115:0] concat_1140;
wire [16:0] add_1329;
wire [19:0] addW_1518;
wire [8:0] slice_1707;
wire [44:0] concat_1896;
wire [22:0] lsl_68;
wire [64:0] subW_257;
wire [13:0] mul_446;
wire [4:0] slice_635;
wire [9:0] mul_824;
wire [11:0] addW_1013;
wire [59:0] concat_1202;
wire [29:0] concat_1391;
wire [7:0] slice_1580;
wire [15:0] lsl_1769;
wire [11:0] addW_1958;
wire [9:0] mul_130;
wire [16:0] add_319;
wire [30:0] concat_508;
wire [112:0] slice_697;
wire [18:0] lsl_886;
wire [58:0] concat_1075;
wire [11:0] slice_1264;
wire [11:0] addW_1453;
wire [4:0] slice_1642;
wire [13:0] mul_1831;
wire [11:0] mul_192;
wire [21:0] concat_381;
wire [6:0] slice_570;
wire [27:0] slice_759;
wire [19:0] addW_948;
wire [61:0] subW_1137;
wire [10:0] add_1326;
wire [35:0] mul_1515;
wire [19:0] add_1704;
wire [6:0] slice_1893;
wire [13:0] mulnw_65;
wire [17:0] slice_254;
wire [13:0] mul_443;
wire [43:0] concat_632;
wire [8:0] mulnw_821;
wire [14:0] concat_1010;
wire [30:0] addW_1199;
wire [15:0] addW_1388;
wire [56:0] slice_1577;
wire [4:0] slice_1766;
wire [14:0] concat_1955;
wire [9:0] mul_127;
wire [10:0] add_316;
wire [16:0] addW_505;
wire [173:0] addW_694;
wire [30:0] concat_883;
wire [42:0] subW_1072;
wire [28:0] slice_1261;
wire [14:0] concat_1450;
wire [4:0] slice_1639;
wire [13:0] mul_1828;
assign slice_189 = mul_188[11:6];
assign addW_378 = mul_376 + mul_377;
assign slice_567 = slice_549[13:0];
assign addW_756 = concat_736 + addW_755;
assign addW_945 = slice_940 + slice_922;
assign slice_1134 = concat_1111[13:0];
assign slice_1323 = slice_1304[4:0];
assign concat_1512 = {addW_1510,slice_1511};
assign lsl_1701 = add_1700 << 5;
assign mul_1890 = slice_1884 * slice_1882;
assign subW_251 = concat_250 - concat_196;
assign slice_440 = slice_439[13:7];
assign slice_629 = addW_613[17:0];
assign lsl_818 = mulnw_817 << 10;
assign slice_1007 = slice_1003[4:0];
assign mul_1196 = slice_1168 * slice_1153;
assign concat_1385 = {mul_1380,slice_1384};
assign addW_1574 = concat_1494 + subW_1573;
assign mulnw_1763 = slice_1741 * slice_1762;
assign slice_1952 = slice_1948[4:0];
assign mul_124 = slice_120 * slice_123;
assign mulnw_313 = slice_294 * slice_310;
assign concat_502 = {mul_497,slice_501};
assign concat_691 = {addW_689,slice_690};
assign slice_880 = addW_864[8:0];
assign slice_1069 = mul_1042[8:0];
assign addW_1258 = concat_1238 + addW_1257;
assign slice_1447 = slice_1443[4:0];
assign concat_1636 = {addW_1634,slice_1635};
assign mul_1825 = slice_1822 * slice_1824;
assign slice_186 = slice_180[5:0];
assign concat_375 = {mul_370,slice_374};
assign addW_564 = concat_560 + addW_563;
assign add_753 = lsl_751 + mul_752;
assign mul_942 = slice_940 * slice_941;
assign add_1131 = lsl_1124 + add_1130;
assign slice_1320 = slice_1304[8:5];
assign addW_1509 = mul_1507 + mul_1508;
assign mulnw_1698 = slice_1697 * slice_1665;
assign slice_1887 = mul_1886[13:7];
assign addW_248 = concat_224 + addW_247;
assign slice_437 = mul_430[6:0];
assign slice_626 = mul_619[5:0];
assign add_815 = lsl_807 + add_814;
assign slice_1004 = slice_1003[9:5];
assign mulnw_1193 = slice_1164 * slice_1153;
assign slice_1382 = slice_1378[6:0];
assign concat_1571 = {addW_1569,slice_1570};
assign slice_1760 = mul_1759[17:9];
assign slice_1949 = slice_1948[9:5];
assign addW_121 = slice_111 + slice_93;
assign slice_310 = slice_306[8:5];
assign slice_499 = slice_495[6:0];
assign subW_688 = subW_687 - concat_606;
assign slice_877 = mul_870[4:0];
assign add_1066 = lsl_1058 + add_1065;
assign add_1255 = lsl_1253 + mul_1254;
assign slice_1444 = slice_1443[9:5];
assign addW_1633 = add_1623 + add_1632;
assign slice_1822 = slice_1821[13:7];
assign slice_2011 = concat_1349[112:0];
assign slice_183 = addW_182[29:18];
assign slice_372 = slice_368[4:0];
assign mul4_561 = slice_551 * slice_557;
assign add_750 = mulnw_748 + mulnw_749;
assign concat_939 = {addW_937,slice_938};
assign lsl_1128 = add_1127 << 7;
assign mul_1317 = slice_1293 * slice_1313;
assign concat_1506 = {mul_1501,slice_1505};
assign mulnw_1695 = slice_1694 * slice_1665;
assign slice_1884 = slice_1879[6:0];
assign addW_56 = concat_51 + addW_55;
assign add_245 = lsl_243 + mul_244;
assign mul4_434 = slice_428 * slice_426;
assign mul_623 = slice_617 * slice_615;
assign lsl_812 = add_811 << 5;
assign slice_1001 = slice_1000[9:5];
assign mulnw_1190 = slice_1164 * slice_1150;
assign slice_1379 = slice_1378[13:7];
assign subW_1568 = subW_1567 - mul_1515;
assign slice_1757 = addW_1739[8:0];
assign slice_1946 = slice_1945[9:5];
assign addW_118 = slice_110 + slice_89;
assign mul_307 = slice_305 * slice_306;
assign slice_496 = slice_495[14:7];
assign slice_685 = mul_630[17:0];
assign mul_874 = slice_868 * slice_866;
assign lsl_1063 = add_1062 << 5;
assign add_1252 = mulnw_1250 + mulnw_1251;
assign slice_1441 = slice_1440[9:5];
assign mul_1630 = slice_1602 * slice_1587;
assign slice_1819 = mul_1812[6:0];
assign subW_2008 = concat_2007 - concat_696;
assign slice_180 = addW_179[29:18];
assign slice_369 = slice_368[9:5];
assign mul_558 = slice_556 * slice_557;
assign lsl_747 = mulnw_746 << 14;
assign addW_936 = mul_934 + mul_935;
assign mulnw_1125 = slice_1101 * slice_1083;
assign mulnw_1314 = slice_1288 * slice_1313;
assign slice_1503 = slice_1499[5:0];
assign add_1692 = lsl_1690 + mul_1691;
assign slice_1881 = slice_1864[13:0];
assign mul_53 = slice_43 * slice_48;
assign add_242 = mulnw_240 + mulnw_241;
assign slice_431 = mul_430[13:7];
assign slice_620 = mul_619[11:6];
assign slice_809 = slice_801[4:0];
assign concat_998 = {addW_996,slice_997};
assign mul_1187 = slice_1152 * slice_1169;
assign slice_1376 = slice_1356[13:0];
assign slice_1565 = mul_1538[8:0];
assign addW_1754 = concat_1750 + addW_1753;
assign concat_1943 = {concat_1938,slice_1942};
assign concat_115 = {concat_108,slice_114};
assign concat_304 = {addW_302,slice_303};
assign addW_493 = slice_266 + slice_21;
assign subW_682 = concat_681 - concat_627;
assign slice_871 = mul_870[9:5];
assign mulnw_1060 = slice_1059 * slice_1027;
assign lsl_1249 = mulnw_1248 << 14;
assign concat_1438 = {concat_1433,slice_1437};
assign mulnw_1627 = slice_1598 * slice_1587;
assign mul4_1816 = slice_1810 * slice_1808;
assign addW_2005 = concat_1799 + subW_2004;
assign slice_366 = slice_365[9:5];
assign mul_555 = slice_551 * slice_554;
assign add_744 = lsl_742 + mul_743;
assign concat_933 = {mul_928,slice_932};
assign add_1122 = lsl_1115 + add_1121;
assign lsl_1311 = mulnw_1310 << 10;
assign slice_1500 = slice_1499[11:6];
assign add_1689 = mulnw_1686 + mulnw_1688;
assign concat_1878 = {addW_1876,slice_1877};
assign slice_50 = mul_49[13:7];
assign slice_239 = slice_220[4:0];
assign slice_428 = slice_422[6:0];
assign slice_617 = slice_611[5:0];
assign mulnw_806 = slice_784 * slice_805;
assign subW_995 = subW_994 - mul_942;
assign mulnw_1184 = slice_1146 * slice_1169;
assign addW_1373 = concat_1369 + addW_1372;
assign add_1562 = lsl_1554 + add_1561;
assign mul_1751 = slice_1741 * slice_1747;
assign slice_1940 = addW_1924[17:0];
assign mul_112 = slice_110 * slice_111;
assign addW_301 = mul_299 + mul_300;
assign slice_490 = addW_489[57:29];
assign addW_679 = concat_655 + addW_678;
assign slice_868 = slice_862[4:0];
assign mulnw_1057 = slice_1056 * slice_1027;
assign add_1246 = lsl_1244 + mul_1245;
assign slice_1435 = slice_1419[17:0];
assign mulnw_1624 = slice_1598 * slice_1584;
assign slice_1813 = mul_1812[13:7];
assign concat_2002 = {addW_2000,slice_2001};
assign concat_363 = {concat_358,slice_362};
assign slice_552 = addW_493[28:0];
assign add_741 = mulnw_739 + mulnw_740;
assign slice_930 = slice_926[4:0];
assign lsl_1119 = add_1118 << 7;
assign concat_1308 = {concat_1303,slice_1307};
assign slice_1497 = slice_1496[11:6];
assign mulnw_1686 = slice_1667 * slice_1683;
assign addW_1875 = mul4_1873 + mul4_1874;
assign slice_47 = slice_42[6:0];
assign slice_236 = slice_220[8:5];
assign slice_425 = addW_424[28:14];
assign slice_614 = addW_613[29:18];
assign slice_803 = mul_802[17:9];
assign slice_992 = mul_965[8:0];
assign mulnw_1181 = slice_1146 * slice_1166;
assign mul4_1370 = slice_1358 * slice_1366;
assign lsl_1559 = add_1558 << 5;
assign mul_1748 = slice_1746 * slice_1747;
assign slice_1937 = mul_1930[5:0];
assign concat_298 = {mul_293,slice_297};
assign add_676 = lsl_674 + mul_675;
assign slice_865 = addW_864[18:9];
assign add_1054 = lsl_1052 + mul_1053;
assign add_1243 = mulnw_1241 + mulnw_1242;
assign slice_1432 = mul_1425[4:0];
assign mul_1621 = slice_1586 * slice_1603;
assign slice_1810 = slice_1803[6:0];
assign subW_1999 = subW_1998 - concat_1918;
assign addW_171 = concat_115 + subW_170;
assign slice_360 = slice_344[17:0];
assign slice_549 = addW_489[28:0];
assign lsl_738 = mulnw_737 << 14;
assign slice_927 = slice_926[9:5];
assign mulnw_1116 = slice_1085 * slice_1099;
assign slice_1305 = addW_1289[8:0];
assign concat_1494 = {concat_1415,slice_1493};
assign slice_1683 = slice_1679[8:5];
assign concat_1872 = {mul_1867,slice_1871};
assign slice_44 = slice_22[13:0];
assign mul_233 = slice_209 * slice_229;
assign slice_422 = addW_421[28:14];
assign slice_611 = addW_610[29:18];
assign slice_800 = addW_782[8:0];
assign add_989 = lsl_981 + add_988;
assign concat_1178 = {addW_1176,slice_1177};
assign mul_1367 = slice_1365 * slice_1366;
assign mulnw_1556 = slice_1555 * slice_1523;
assign mul_1745 = slice_1741 * slice_1744;
assign mul_1934 = slice_1928 * slice_1926;
assign addW_106 = concat_101 + addW_105;
assign slice_295 = slice_291[4:0];
assign add_673 = mulnw_671 + mulnw_672;
assign slice_862 = addW_861[18:9];
assign add_1051 = mulnw_1048 + mulnw_1050;
assign lsl_1240 = mulnw_1239 << 14;
assign mul_1429 = slice_1423 * slice_1421;
assign mulnw_1618 = slice_1580 * slice_1603;
assign slice_1807 = slice_1806[28:14];
assign slice_1996 = mul_1941[17:0];
assign concat_168 = {addW_166,slice_167};
assign slice_357 = mul_350[4:0];
assign addW_546 = concat_526 + addW_545;
assign slice_735 = concat_734[27:14];
assign slice_924 = slice_702[55:0];
assign concat_1113 = {concat_1095,slice_1112};
assign slice_1302 = mul_1295[4:0];
assign slice_1491 = mul_1436[17:0];
assign mul_1680 = slice_1678 * slice_1679;
assign slice_1869 = slice_1865[6:0];
assign mulnw_230 = slice_204 * slice_229;
assign concat_419 = {concat_340,slice_418};
assign concat_608 = {concat_548,slice_607};
assign addW_797 = concat_793 + addW_796;
assign lsl_986 = add_985 << 5;
assign addW_1175 = mul_1173 + mul_1174;
assign mul_1364 = slice_1358 * slice_1363;
assign mulnw_1553 = slice_1552 * slice_1523;
assign addW_1742 = slice_1735 + slice_1720;
assign slice_1931 = mul_1930[11:6];
assign mul_103 = slice_91 * slice_98;
assign slice_292 = slice_291[9:5];
assign addW_481 = concat_419 + subW_480;
assign slice_670 = slice_651[4:0];
assign slice_859 = mul_858[35:18];
assign mulnw_1048 = slice_1029 * slice_1045;
assign slice_1237 = concat_1236[27:14];
assign slice_1426 = mul_1425[9:5];
assign mulnw_1615 = slice_1580 * slice_1600;
assign slice_1804 = slice_1803[14:7];
assign subW_1993 = concat_1992 - concat_1938;
assign addW_165 = add_153 + add_164;
assign mul_354 = slice_348 * slice_346;
assign add_543 = lsl_541 + mul_542;
assign addW_732 = concat_728 + addW_731;
assign slice_921 = slice_920[55:28];
assign slice_1110 = mul_1103[6:0];
assign mul_1299 = slice_1293 * slice_1291;
assign subW_1488 = concat_1487 - concat_1433;
assign concat_1677 = {addW_1675,slice_1676};
assign slice_1866 = slice_1865[14:7];
assign addW_38 = concat_33 + addW_37;
assign lsl_227 = mulnw_226 << 10;
assign slice_416 = mul_361[17:0];
assign slice_605 = concat_582[13:0];
assign mul_794 = slice_784 * slice_790;
assign mulnw_983 = slice_982 * slice_950;
assign concat_1172 = {mul_1167,slice_1171};
assign slice_1361 = slice_1360[56:28];
assign add_1550 = lsl_1548 + mul_1549;
assign addW_1739 = slice_1734 + slice_1717;
assign slice_1928 = slice_1922[5:0];
assign slice_100 = mul_99[9:5];
assign slice_289 = slice_288[9:5];
assign concat_478 = {addW_476,slice_477};
assign slice_667 = slice_651[8:5];
assign slice_856 = addW_838[17:0];
assign slice_1045 = slice_1041[8:5];
assign addW_1234 = concat_1230 + addW_1233;
assign slice_1423 = slice_1417[4:0];
assign concat_1612 = {addW_1610,slice_1611};
assign addW_1801 = slice_1577 + slice_1355;
assign addW_1990 = concat_1966 + addW_1989;
assign mul_162 = slice_157 * slice_126;
assign slice_351 = mul_350[9:5];
assign add_540 = mulnw_538 + mulnw_539;
assign mul_729 = slice_720 * slice_725;
assign slice_918 = concat_835[27:0];
assign mul_1107 = slice_1101 * slice_1099;
assign slice_1296 = mul_1295[9:5];
assign addW_1485 = concat_1461 + addW_1484;
assign addW_1674 = mul_1672 + mul_1673;
assign slice_1863 = slice_1862[14:7];
assign mul4_35 = slice_18 * slice_29;
assign concat_224 = {concat_219,slice_223};
assign subW_413 = concat_412 - concat_358;
assign add_602 = lsl_595 + add_601;
assign mul_791 = slice_789 * slice_790;
assign mulnw_980 = slice_979 * slice_950;
assign slice_1169 = slice_1165[6:0];
assign slice_1358 = slice_1357[14:7];
assign add_1547 = mulnw_1544 + mulnw_1546;
assign mul_1736 = slice_1734 * slice_1735;
assign slice_1925 = addW_1924[29:18];
assign slice_97 = slice_89[4:0];
assign concat_286 = {concat_281,slice_285};
assign addW_475 = add_465 + add_474;
assign mul_664 = slice_640 * slice_660;
assign addW_853 = concat_849 + addW_852;
assign mul_1042 = slice_1040 * slice_1041;
assign mul_1231 = slice_1222 * slice_1227;
assign slice_1420 = slice_1419[27:18];
assign addW_1609 = mul_1607 + mul_1608;
assign slice_1798 = concat_1797[113:57];
assign add_1987 = lsl_1985 + mul_1986;
assign mulnw_159 = slice_154 * slice_126;
assign slice_348 = slice_342[4:0];
assign lsl_537 = mulnw_536 << 14;
assign mul_726 = slice_724 * slice_725;
assign subW_915 = concat_914 - concat_758;
assign slice_1104 = mul_1103[13:7];
assign slice_1293 = slice_1287[4:0];
assign add_1482 = lsl_1480 + mul_1481;
assign concat_1671 = {mul_1666,slice_1670};
assign concat_1860 = {addW_1858,slice_1859};
assign slice_32 = mul_30[13:7];
assign slice_221 = addW_205[8:0];
assign addW_410 = concat_386 + addW_409;
assign lsl_599 = add_598 << 7;
assign mul_788 = slice_784 * slice_787;
assign add_977 = lsl_975 + mul_976;
assign slice_1166 = slice_1165[13:7];
assign slice_1355 = addW_1354[113:57];
assign mulnw_1544 = slice_1525 * slice_1541;
assign concat_1733 = {addW_1731,slice_1732};
assign slice_1922 = addW_1921[29:18];
assign slice_94 = slice_93[9:5];
assign slice_283 = slice_267[17:0];
assign mul_472 = slice_444 * slice_429;
assign mulnw_661 = slice_635 * slice_660;
assign mul_850 = slice_840 * slice_846;
assign concat_1039 = {addW_1037,slice_1038};
assign mul_1228 = slice_1226 * slice_1227;
assign slice_1417 = slice_1416[27:18];
assign concat_1606 = {mul_1601,slice_1605};
assign addW_1795 = concat_1715 + subW_1794;
assign add_1984 = mulnw_1982 + mulnw_1983;
assign lsl_156 = mulnw_155 << 10;
assign slice_345 = slice_344[27:18];
assign add_534 = lsl_532 + mul_533;
assign mul_723 = slice_720 * slice_722;
assign addW_912 = concat_860 + subW_911;
assign slice_1101 = slice_1096[6:0];
assign slice_1290 = addW_1289[18:9];
assign add_1479 = mulnw_1477 + mulnw_1478;
assign slice_1668 = slice_1664[4:0];
assign addW_1857 = add_1847 + add_1856;
assign slice_29 = slice_23[6:0];
assign slice_218 = mul_211[4:0];
assign add_407 = lsl_405 + mul_406;
assign mulnw_596 = slice_572 * slice_554;
assign addW_785 = slice_778 + slice_763;
assign add_974 = mulnw_971 + mulnw_973;
assign slice_1163 = slice_1144[13:0];
assign slice_1541 = slice_1537[8:5];
assign addW_1730 = mul_1728 + mul_1729;
assign slice_1919 = concat_1918[57:29];
assign slice_91 = slice_89[9:5];
assign slice_280 = mul_273[4:0];
assign mulnw_469 = slice_440 * slice_429;
assign lsl_658 = mulnw_657 << 10;
assign mul_847 = slice_845 * slice_846;
assign addW_1036 = mul_1034 + mul_1035;
assign mul_1225 = slice_1222 * slice_1224;
assign slice_1414 = concat_1391[13:0];
assign slice_1603 = slice_1599[6:0];
assign concat_1792 = {addW_1790,slice_1791};
assign slice_1981 = slice_1962[4:0];
assign add_153 = lsl_145 + add_152;
assign slice_342 = slice_341[27:18];
assign add_531 = mulnw_529 + mulnw_530;
assign slice_720 = slice_719[13:7];
assign concat_909 = {addW_907,slice_908};
assign slice_1098 = addW_1081[13:0];
assign slice_1287 = addW_1286[18:9];
assign slice_1476 = slice_1457[4:0];
assign slice_1665 = slice_1664[9:5];
assign mul_1854 = slice_1826 * slice_1811;
assign mul_215 = slice_209 * slice_207;
assign add_404 = mulnw_402 + mulnw_403;
assign add_593 = lsl_586 + add_592;
assign addW_782 = slice_777 + slice_760;
assign mulnw_971 = slice_952 * slice_968;
assign addW_1160 = concat_1156 + addW_1159;
assign concat_1349 = {addW_1347,slice_1348};
assign mul_1538 = slice_1536 * slice_1537;
assign concat_1727 = {mul_1722,slice_1726};
assign addW_1916 = concat_1896 + addW_1915;
assign mul_277 = slice_271 * slice_269;
assign mulnw_466 = slice_440 * slice_426;
assign concat_655 = {concat_650,slice_654};
assign mul_844 = slice_840 * slice_843;
assign concat_1033 = {mul_1028,slice_1032};
assign slice_1222 = slice_1221[13:7];
assign add_1411 = lsl_1404 + add_1410;
assign slice_1600 = slice_1599[13:7];
assign subW_1789 = subW_1788 - mul_1736;
assign slice_1978 = slice_1962[8:5];
assign lsl_150 = add_149 << 5;
assign slice_339 = mul_284[17:0];
assign lsl_528 = mulnw_527 << 14;
assign slice_717 = mul_710[6:0];
assign addW_906 = add_894 + add_905;
assign concat_1095 = {addW_1093,slice_1094};
assign slice_1284 = mul_1283[35:18];
assign slice_1473 = slice_1457[8:5];
assign slice_1662 = slice_1661[9:5];
assign mulnw_1851 = slice_1822 * slice_1811;
assign slice_23 = slice_22[28:14];
assign slice_212 = mul_211[9:5];
assign slice_401 = slice_382[4:0];
assign lsl_590 = add_589 << 7;
assign mul_779 = slice_777 * slice_778;
assign slice_968 = slice_964[8:5];
assign mul4_1157 = slice_1146 * slice_1153;
assign subW_1346 = subW_1345 - concat_1140;
assign concat_1535 = {addW_1533,slice_1534};
assign slice_1724 = slice_1720[5:0];
assign add_1913 = lsl_1911 + mul_1912;
assign slice_274 = mul_273[9:5];
assign mul_463 = slice_428 * slice_445;
assign slice_652 = addW_636[8:0];
assign addW_841 = slice_762 + slice_704;
assign slice_1030 = slice_1026[4:0];
assign slice_1219 = mul_1212[6:0];
assign lsl_1408 = add_1407 << 7;
assign slice_1597 = slice_1578[13:0];
assign slice_1786 = mul_1759[8:0];
assign mul_1975 = slice_1951 * slice_1971;
assign slice_147 = slice_137[4:0];
assign subW_336 = concat_335 - concat_281;
assign slice_525 = concat_524[27:14];
assign mul4_714 = slice_708 * slice_706;
assign mul_903 = slice_898 * slice_869;
assign addW_1092 = mul4_1090 + mul4_1091;
assign slice_1281 = addW_1263[17:0];
assign mul_1470 = slice_1446 * slice_1466;
assign concat_1659 = {concat_1654,slice_1658};
assign mulnw_1848 = slice_1822 * slice_1808;
assign slice_20 = IN2[225:113];
assign slice_209 = slice_203[4:0];
assign slice_398 = slice_382[8:5];
assign mulnw_587 = slice_556 * slice_570;
assign concat_776 = {addW_774,slice_775};
assign mul_965 = slice_963 * slice_964;
assign mul_1154 = slice_1152 * slice_1153;
assign slice_1343 = concat_1260[28:0];
assign addW_1532 = mul_1530 + mul_1531;
assign slice_1721 = slice_1720[11:6];
assign add_1910 = mulnw_1908 + mulnw_1909;
assign addW_82 = concat_61 + addW_81;
assign slice_271 = slice_264[4:0];
assign mulnw_460 = slice_423 * slice_445;
assign slice_649 = mul_642[4:0];
assign addW_838 = slice_759 + slice_699;
assign slice_1027 = slice_1026[9:5];
assign mul4_1216 = slice_1210 * slice_1208;
assign mulnw_1405 = slice_1381 * slice_1363;
assign addW_1594 = concat_1590 + addW_1593;
assign add_1783 = lsl_1775 + add_1782;
assign mulnw_1972 = slice_1946 * slice_1971;
assign mulnw_144 = slice_120 * slice_143;
assign addW_333 = concat_309 + addW_332;
assign addW_522 = concat_518 + addW_521;
assign slice_711 = mul_710[13:7];
assign mulnw_900 = slice_895 * slice_869;
assign concat_1089 = {mul_1084,slice_1088};
assign addW_1278 = concat_1274 + addW_1277;
assign mulnw_1467 = slice_1441 * slice_1466;
assign slice_1656 = slice_1640[17:0];
assign mul_1845 = slice_1810 * slice_1827;
assign slice_206 = addW_205[18:9];
assign mul_395 = slice_371 * slice_391;
assign concat_584 = {concat_566,slice_583};
assign addW_773 = mul_771 + mul_772;
assign concat_962 = {addW_960,slice_961};
assign mul_1151 = slice_1146 * slice_1150;
assign subW_1340 = concat_1339 - concat_1202;
assign concat_1529 = {mul_1524,slice_1528};
assign slice_1718 = slice_1717[11:6];
assign lsl_1907 = mulnw_1906 << 14;
assign add_79 = lsl_77 + mul_78;
assign slice_268 = slice_267[27:18];
assign mulnw_457 = slice_423 * slice_442;
assign mul_646 = slice_640 * slice_638;
assign concat_835 = {addW_833,slice_834};
assign slice_1024 = slice_1023[9:5];
assign slice_1213 = mul_1212[13:7];
assign add_1402 = lsl_1395 + add_1401;
assign mul4_1591 = slice_1580 * slice_1587;
assign lsl_1780 = add_1779 << 5;
assign lsl_1969 = mulnw_1968 << 10;
assign add_330 = lsl_328 + mul_329;
assign mul_519 = slice_510 * slice_515;
assign slice_708 = slice_700[6:0];
assign lsl_897 = mulnw_896 << 10;
assign slice_1086 = slice_1082[6:0];
assign mul_1275 = slice_1265 * slice_1271;
assign lsl_1464 = mulnw_1463 << 10;
assign slice_1653 = mul_1646[4:0];
assign mulnw_1842 = slice_1804 * slice_1827;
assign slice_14 = slice_12[56:28];
assign slice_203 = addW_202[18:9];
assign mulnw_392 = slice_366 * slice_391;
assign slice_581 = mul_574[6:0];
assign concat_770 = {mul_765,slice_769};
assign addW_959 = mul_957 + mul_958;
assign slice_1148 = addW_1147[57:29];
assign addW_1337 = concat_1285 + subW_1336;
assign slice_1526 = slice_1522[4:0];
assign concat_1715 = {concat_1636,slice_1714};
assign add_1904 = lsl_1902 + mul_1903;
assign add_76 = mulnw_74 + mulnw_75;
assign slice_265 = slice_264[9:5];
assign concat_454 = {addW_452,slice_453};
assign slice_643 = mul_642[9:5];
assign subW_832 = subW_831 - mul_779;
assign concat_1021 = {concat_1016,slice_1020};
assign slice_1210 = slice_1204[6:0];
assign lsl_1399 = add_1398 << 7;
assign mul_1588 = slice_1586 * slice_1587;
assign mulnw_1777 = slice_1776 * slice_1744;
assign concat_1966 = {concat_1961,slice_1965};
assign mul_138 = slice_136 * slice_137;
assign add_327 = mulnw_325 + mulnw_326;
assign mul_516 = slice_514 * slice_515;
assign slice_705 = slice_704[28:14];
assign add_894 = lsl_886 + add_893;
assign slice_1083 = slice_1082[14:7];
assign mul_1272 = slice_1270 * slice_1271;
assign concat_1461 = {concat_1456,slice_1460};
assign mul_1650 = slice_1644 * slice_1642;
assign mulnw_1839 = slice_1804 * slice_1824;
assign slice_200 = mul_199[35:18];
assign lsl_389 = mulnw_388 << 10;
assign mul_578 = slice_572 * slice_570;
assign slice_767 = slice_763[4:0];
assign concat_956 = {mul_951,slice_955};
assign slice_1145 = slice_1144[28:14];
assign concat_1334 = {addW_1332,slice_1333};
assign slice_1523 = slice_1522[9:5];
assign slice_1712 = mul_1657[17:0];
assign add_1901 = mulnw_1899 + mulnw_1900;
assign lsl_73 = mulnw_72 << 14;
assign slice_262 = slice_9[55:0];
assign addW_451 = mul_449 + mul_450;
assign slice_640 = slice_634[4:0];
assign slice_829 = mul_802[8:0];
assign slice_1018 = slice_1002[17:0];
assign slice_1207 = slice_1206[28:14];
assign mulnw_1396 = slice_1365 * slice_1379;
assign mul_1585 = slice_1580 * slice_1584;
assign mulnw_1774 = slice_1773 * slice_1744;
assign slice_1963 = addW_1947[8:0];
assign concat_135 = {addW_133,slice_134};
assign slice_324 = slice_305[4:0];
assign mul_513 = slice_510 * slice_512;
assign slice_702 = IN2[112:0];
assign lsl_891 = add_890 << 5;
assign slice_1080 = slice_1079[14:7];
assign mul_1269 = slice_1265 * slice_1268;
assign slice_1458 = addW_1442[8:0];
assign slice_1647 = mul_1646[9:5];
assign concat_1836 = {addW_1834,slice_1835};
assign slice_197 = addW_179[17:0];
assign concat_386 = {concat_381,slice_385};
assign slice_575 = mul_574[13:7];
assign slice_764 = slice_763[9:5];
assign slice_953 = slice_949[4:0];
assign concat_1142 = {concat_919,slice_1141};
assign addW_1331 = add_1319 + add_1330;
assign slice_1520 = slice_1519[9:5];
assign subW_1709 = concat_1708 - concat_1654;
assign lsl_1898 = mulnw_1897 << 14;
assign add_70 = lsl_68 + mul_69;
assign slice_259 = concat_173[27:0];
assign concat_448 = {mul_443,slice_447};
assign slice_637 = addW_636[18:9];
assign add_826 = lsl_818 + add_825;
assign slice_1015 = mul_1008[4:0];
assign slice_1204 = slice_1203[28:14];
assign concat_1393 = {concat_1375,slice_1392};
assign slice_1582 = slice_1581[56:28];
assign add_1771 = lsl_1769 + mul_1770;
assign slice_1960 = mul_1953[4:0];
assign addW_132 = mul_130 + mul_131;
assign slice_321 = slice_305[8:5];
assign slice_510 = slice_509[13:7];
assign slice_699 = slice_698[56:28];
assign slice_888 = slice_880[4:0];
assign concat_1077 = {concat_998,slice_1076};
assign addW_1266 = slice_1206 + slice_1148;
assign slice_1455 = mul_1448[4:0];
assign slice_1644 = slice_1638[4:0];
assign addW_1833 = mul_1831 + mul_1832;
assign addW_194 = concat_190 + addW_193;
assign slice_383 = addW_367[8:0];
assign slice_572 = slice_567[6:0];
assign slice_761 = slice_760[9:5];
assign slice_950 = slice_949[9:5];
assign slice_1139 = concat_1075[27:0];
assign mul_1328 = slice_1323 * slice_1294;
assign concat_1517 = {concat_1512,slice_1516};
assign addW_1706 = concat_1682 + addW_1705;
assign slice_1895 = concat_1894[27:14];
assign add_67 = mulnw_65 + mulnw_66;
assign subW_256 = concat_255 - concat_84;
assign slice_445 = slice_441[6:0];
assign slice_634 = addW_633[18:9];
assign lsl_823 = add_822 << 5;
assign mul_1012 = slice_1006 * slice_1004;
assign slice_1201 = concat_1178[13:0];
assign slice_1390 = mul_1383[6:0];
assign slice_1579 = slice_1578[28:14];
assign add_1768 = mulnw_1765 + mulnw_1767;
assign mul_1957 = slice_1951 * slice_1949;
assign concat_129 = {mul_124,slice_128};
assign mul_318 = slice_294 * slice_314;
assign slice_507 = mul_500[6:0];
assign concat_696 = {addW_694,slice_695};
assign mulnw_885 = slice_863 * slice_884;
assign slice_1074 = mul_1019[17:0];
assign addW_1263 = slice_1203 + slice_1144;
assign mul_1452 = slice_1446 * slice_1444;
assign slice_1641 = slice_1640[27:18];
assign concat_1830 = {mul_1825,slice_1829};
assign mul_191 = slice_181 * slice_187;
assign slice_380 = mul_373[4:0];
assign slice_569 = slice_552[13:0];
assign concat_758 = {addW_756,slice_757};
assign slice_947 = slice_946[9:5];
assign subW_1136 = concat_1135 - concat_998;
assign mulnw_1325 = slice_1320 * slice_1294;
assign slice_1514 = addW_1498[17:0];
assign add_1703 = lsl_1701 + mul_1702;
assign addW_1892 = concat_1888 + addW_1891;
assign lsl_64 = mulnw_63 << 14;
assign addW_253 = concat_201 + subW_252;
assign slice_442 = slice_441[13:7];
assign slice_631 = mul_630[35:18];
assign mulnw_820 = slice_819 * slice_787;
assign slice_1009 = mul_1008[9:5];
assign add_1198 = lsl_1191 + add_1197;
assign mul_1387 = slice_1381 * slice_1379;
assign concat_1576 = {addW_1574,slice_1575};
assign mulnw_1765 = slice_1746 * slice_1762;
assign slice_1954 = mul_1953[9:5];
assign slice_126 = slice_122[4:0];
assign mulnw_315 = slice_289 * slice_314;
assign mul4_504 = slice_498 * slice_496;
assign subW_693 = subW_692 - concat_483;
assign slice_882 = mul_881[17:9];
assign subW_1071 = concat_1070 - concat_1016;
assign concat_1260 = {addW_1258,slice_1259};
assign slice_1449 = mul_1448[9:5];
assign slice_1638 = slice_1637[27:18];
assign slice_1827 = slice_1823[6:0];
assign mul_188 = slice_186 * slice_187;
assign mul_377 = slice_371 * slice_369;
assign concat_566 = {addW_564,slice_565};
assign addW_755 = add_745 + add_754;
assign concat_944 = {concat_939,slice_943};
assign addW_1133 = concat_1113 + addW_1132;
assign lsl_1322 = mulnw_1321 << 10;
assign slice_1511 = mul_1504[5:0];
assign add_1700 = mulnw_1698 + mulnw_1699;
assign mul_1889 = slice_1880 * slice_1885;
assign concat_61 = {concat_40,slice_60};
assign concat_250 = {addW_248,slice_249};
assign slice_439 = addW_421[13:0];
assign slice_628 = addW_610[17:0];
assign mulnw_817 = slice_816 * slice_787;
assign slice_1006 = slice_1000[4:0];
assign lsl_1195 = add_1194 << 7;
assign slice_1384 = mul_1383[13:7];
assign subW_1573 = subW_1572 - concat_1492;
assign slice_1762 = slice_1758[8:5];
assign slice_1951 = slice_1945[4:0];
assign slice_123 = slice_122[9:5];
assign lsl_312 = mulnw_311 << 10;
assign slice_501 = mul_500[13:7];
assign slice_690 = concat_606[28:0];
assign slice_879 = addW_861[8:0];
assign addW_1068 = concat_1044 + addW_1067;
assign addW_1257 = add_1247 + add_1256;
assign slice_1446 = slice_1440[4:0];
assign slice_1635 = concat_1612[13:0];
assign slice_1824 = slice_1823[13:7];
assign mul_185 = slice_181 * slice_184;
assign slice_374 = mul_373[9:5];
assign addW_563 = mul4_561 + mul4_562;
assign mul_752 = slice_724 * slice_709;
assign slice_941 = slice_925[17:0];
assign add_1130 = lsl_1128 + mul_1129;
assign add_1319 = lsl_1311 + add_1318;
assign mul_1508 = slice_1502 * slice_1500;
assign slice_1697 = slice_1678[4:0];
assign mul_1886 = slice_1884 * slice_1885;
assign concat_58 = {addW_56,slice_57};
assign addW_247 = add_235 + add_246;
assign addW_436 = concat_432 + addW_435;
assign addW_625 = concat_621 + addW_624;
assign add_814 = lsl_812 + mul_813;
assign slice_1003 = slice_1002[27:18];
assign mulnw_1192 = slice_1168 * slice_1150;
assign slice_1381 = slice_1376[6:0];
assign slice_1570 = mul_1515[17:0];
assign mul_1759 = slice_1757 * slice_1758;
assign slice_1948 = addW_1947[18:9];
assign slice_120 = slice_119[9:5];
assign concat_309 = {concat_304,slice_308};
assign slice_498 = slice_491[6:0];
assign subW_687 = concat_686 - concat_548;
assign addW_876 = concat_872 + addW_875;
assign add_1065 = lsl_1063 + mul_1064;
assign mul_1254 = slice_1226 * slice_1211;
assign slice_1443 = addW_1442[18:9];
assign add_1632 = lsl_1625 + add_1631;
assign slice_1821 = slice_1802[13:0];
assign addW_2010 = concat_1351 + subW_2009;
assign addW_182 = slice_92 + slice_22;
assign slice_371 = slice_365[4:0];
assign concat_560 = {mul_555,slice_559};
assign mulnw_749 = slice_720 * slice_709;
assign slice_938 = mul_931[4:0];
assign add_1127 = mulnw_1125 + mulnw_1126;
assign lsl_1316 = add_1315 << 5;
assign slice_1505 = mul_1504[11:6];
assign slice_1694 = slice_1678[8:5];
assign mul_1883 = slice_1880 * slice_1882;
assign addW_55 = mul_53 + mul_54;
assign mul_244 = slice_239 * slice_210;
assign mul4_433 = slice_423 * slice_429;
assign mul_622 = slice_612 * slice_618;
assign add_811 = mulnw_808 + mulnw_810;
assign slice_1000 = slice_999[27:18];
assign add_1189 = lsl_1182 + add_1188;
assign slice_1378 = slice_1361[13:0];
assign subW_1567 = concat_1566 - concat_1512;
assign concat_1756 = {addW_1754,slice_1755};
assign slice_1945 = addW_1944[18:9];
assign slice_306 = addW_290[8:0];
assign slice_495 = slice_494[28:14];
assign addW_684 = concat_632 + subW_683;
assign mul_873 = slice_863 * slice_869;
assign add_1062 = mulnw_1060 + mulnw_1061;
assign mulnw_1251 = slice_1222 * slice_1211;
assign slice_1440 = addW_1439[18:9];
assign lsl_1629 = add_1628 << 7;
assign addW_1818 = concat_1814 + addW_1817;
assign concat_2007 = {addW_2005,slice_2006};
assign addW_179 = slice_87 + slice_14;
assign slice_368 = addW_367[18:9];
assign slice_557 = slice_553[6:0];
assign mulnw_746 = slice_720 * slice_706;
assign mul_935 = slice_929 * slice_927;
assign lsl_1124 = mulnw_1123 << 14;
assign slice_1313 = slice_1305[4:0];
assign slice_1502 = slice_1496[5:0];
assign mul_1691 = slice_1667 * slice_1687;
assign slice_1880 = slice_1879[13:7];
assign mulnw_241 = slice_236 * slice_210;
assign mul_430 = slice_428 * slice_429;
assign mul_619 = slice_617 * slice_618;
assign mulnw_808 = slice_789 * slice_805;
assign slice_997 = mul_942[17:0];
assign lsl_1186 = add_1185 << 7;
assign concat_1375 = {addW_1373,slice_1374};
assign addW_1564 = concat_1540 + addW_1563;
assign addW_1753 = mul_1751 + mul_1752;
assign slice_1942 = mul_1941[35:18];
assign slice_114 = mul_112[35:18];
assign slice_303 = mul_296[4:0];
assign slice_492 = slice_491[14:7];
assign concat_681 = {addW_679,slice_680};
assign mul_870 = slice_868 * slice_869;
assign slice_1059 = slice_1040[4:0];
assign mulnw_1248 = slice_1222 * slice_1208;
assign slice_1437 = mul_1436[35:18];
assign mulnw_1626 = slice_1602 * slice_1584;
assign mul4_1815 = slice_1804 * slice_1811;
assign subW_2004 = subW_2003 - concat_1797;
assign concat_176 = {concat_84,slice_175};
assign slice_365 = addW_364[18:9];
assign slice_554 = slice_553[14:7];
assign mul_743 = slice_708 * slice_725;
assign slice_932 = mul_931[9:5];
assign add_1121 = lsl_1119 + mul_1120;
assign mulnw_1310 = slice_1288 * slice_1309;
assign slice_1499 = addW_1498[29:18];
assign mulnw_1688 = slice_1662 * slice_1687;
assign slice_1877 = mul_1870[6:0];
assign mul_49 = slice_47 * slice_48;
assign lsl_238 = mulnw_237 << 10;
assign mul_427 = slice_423 * slice_426;
assign mul_616 = slice_612 * slice_615;
assign slice_805 = slice_801[8:5];
assign subW_994 = concat_993 - concat_939;
assign mulnw_1183 = slice_1152 * slice_1166;
assign addW_1372 = mul4_1370 + mul4_1371;
assign add_1561 = lsl_1559 + mul_1560;
assign concat_1750 = {mul_1745,slice_1749};
assign slice_1939 = addW_1921[17:0];
assign slice_111 = slice_92[17:0];
assign mul_300 = slice_294 * slice_292;
assign addW_489 = slice_262 + slice_12;
assign addW_678 = add_666 + add_677;
assign mul_867 = slice_863 * slice_866;
assign slice_1056 = slice_1040[8:5];
assign mul_1245 = slice_1210 * slice_1227;
assign slice_1434 = slice_1416[17:0];
assign add_1623 = lsl_1616 + add_1622;
assign mul_1812 = slice_1810 * slice_1811;
assign slice_2001 = concat_1918[28:0];
assign concat_173 = {addW_171,slice_172};
assign slice_362 = mul_361[35:18];
assign slice_551 = slice_550[14:7];
assign mulnw_740 = slice_701 * slice_725;
assign slice_929 = slice_922[4:0];
assign add_1118 = mulnw_1116 + mulnw_1117;
assign slice_1307 = mul_1306[17:9];
assign slice_1496 = addW_1495[29:18];
assign lsl_1685 = mulnw_1684 << 10;
assign mul4_1874 = slice_1868 * slice_1866;
assign mul_46 = slice_43 * slice_45;
assign add_235 = lsl_227 + add_234;
assign addW_424 = slice_344 + slice_267;
assign addW_613 = slice_552 + slice_494;
assign mul_802 = slice_800 * slice_801;
assign addW_991 = concat_967 + addW_990;
assign concat_1180 = {concat_1162,slice_1179};
assign concat_1369 = {mul_1364,slice_1368};
assign add_1558 = mulnw_1556 + mulnw_1557;
assign slice_1747 = slice_1743[4:0];
assign addW_1936 = concat_1932 + addW_1935;
assign concat_108 = {addW_106,slice_107};
assign slice_297 = mul_296[9:5];
assign concat_486 = {concat_260,slice_485};
assign mul_675 = slice_670 * slice_641;
assign addW_864 = slice_857 + slice_842;
assign mul_1053 = slice_1029 * slice_1049;
assign mulnw_1242 = slice_1205 * slice_1227;
assign addW_1431 = concat_1427 + addW_1430;
assign lsl_1620 = add_1619 << 7;
assign mul_1809 = slice_1804 * slice_1808;
assign subW_1998 = concat_1997 - concat_1860;
assign subW_170 = subW_169 - mul_112;
assign slice_359 = slice_341[17:0];
assign concat_548 = {addW_546,slice_547};
assign mulnw_737 = slice_701 * slice_722;
assign slice_926 = slice_925[27:18];
assign lsl_1115 = mulnw_1114 << 14;
assign slice_1304 = addW_1286[8:0];
assign slice_1493 = concat_1492[55:28];
assign concat_1682 = {concat_1677,slice_1681};
assign slice_1871 = mul_1870[13:7];
assign slice_43 = slice_42[13:7];
assign lsl_232 = add_231 << 5;
assign addW_421 = slice_341 + slice_263;
assign addW_610 = slice_549 + slice_490;
assign concat_799 = {addW_797,slice_798};
assign add_988 = lsl_986 + mul_987;
assign slice_1177 = mul_1170[6:0];
assign slice_1366 = slice_1362[6:0];
assign slice_1555 = slice_1536[4:0];
assign slice_1744 = slice_1743[9:5];
assign mul_1933 = slice_1923 * slice_1929;
assign addW_105 = mul_103 + mul_104;
assign slice_294 = slice_288[4:0];
assign concat_483 = {addW_481,slice_482};
assign mulnw_672 = slice_667 * slice_641;
assign addW_861 = slice_856 + slice_839;
assign mulnw_1050 = slice_1024 * slice_1049;
assign mulnw_1239 = slice_1205 * slice_1224;
assign mul_1428 = slice_1418 * slice_1424;
assign mulnw_1617 = slice_1586 * slice_1600;
assign slice_1806 = addW_1805[57:29];
assign addW_1995 = concat_1943 + subW_1994;
assign slice_167 = mul_138[8:0];
assign addW_356 = concat_352 + addW_355;
assign addW_545 = add_535 + add_544;
assign concat_734 = {addW_732,slice_733};
assign slice_923 = slice_922[9:5];
assign slice_1112 = concat_1111[27:14];
assign addW_1301 = concat_1297 + addW_1300;
assign addW_1490 = concat_1438 + subW_1489;
assign slice_1679 = addW_1663[8:0];
assign slice_1868 = slice_1862[6:0];
assign concat_40 = {addW_38,slice_39};
assign slice_229 = slice_221[4:0];
assign slice_418 = concat_417[55:28];
assign slice_607 = concat_606[57:29];
assign addW_796 = mul_794 + mul_795;
assign add_985 = mulnw_983 + mulnw_984;
assign mul_1174 = slice_1168 * slice_1166;
assign slice_1363 = slice_1362[14:7];
assign slice_1552 = slice_1536[8:5];
assign slice_1741 = slice_1740[9:5];
assign mul_1930 = slice_1928 * slice_1929;
assign slice_291 = addW_290[18:9];
assign subW_480 = subW_479 - concat_417;
assign lsl_669 = mulnw_668 << 10;
assign mul_858 = slice_856 * slice_857;
assign lsl_1047 = mulnw_1046 << 10;
assign concat_1236 = {addW_1234,slice_1235};
assign mul_1425 = slice_1423 * slice_1424;
assign concat_1614 = {concat_1596,slice_1613};
assign slice_1803 = slice_1802[28:14];
assign concat_1992 = {addW_1990,slice_1991};
assign add_164 = lsl_156 + add_163;
assign mul_353 = slice_343 * slice_349;
assign mul_542 = slice_514 * slice_499;
assign addW_731 = mul_729 + mul_730;
assign slice_920 = slice_697[55:0];
assign addW_1109 = concat_1105 + addW_1108;
assign mul_1298 = slice_1288 * slice_1294;
assign concat_1487 = {addW_1485,slice_1486};
assign slice_1676 = mul_1669[4:0];
assign slice_1865 = slice_1864[28:14];
assign addW_37 = mul4_35 + mul4_36;
assign mulnw_226 = slice_204 * slice_225;
assign addW_415 = concat_363 + subW_414;
assign addW_604 = concat_584 + addW_603;
assign concat_793 = {mul_788,slice_792};
assign slice_982 = slice_963[4:0];
assign slice_1171 = mul_1170[13:7];
assign slice_1360 = addW_1359[113:57];
assign mul_1549 = slice_1525 * slice_1545;
assign concat_1738 = {concat_1733,slice_1737};
assign mul_1927 = slice_1923 * slice_1926;
assign mul_99 = slice_97 * slice_98;
assign slice_288 = addW_287[18:9];
assign slice_477 = concat_454[13:0];
assign add_666 = lsl_658 + add_665;
assign concat_855 = {addW_853,slice_854};
assign concat_1044 = {concat_1039,slice_1043};
assign addW_1233 = mul_1231 + mul_1232;
assign mul_1422 = slice_1418 * slice_1421;
assign slice_1611 = mul_1604[6:0];
assign addW_1989 = add_1977 + add_1988;
assign lsl_161 = add_160 << 5;
assign mul_350 = slice_348 * slice_349;
assign mulnw_539 = slice_510 * slice_499;
assign concat_728 = {mul_723,slice_727};
assign addW_917 = concat_837 + subW_916;
assign mul_1106 = slice_1097 * slice_1102;
assign mul_1295 = slice_1293 * slice_1294;
assign addW_1484 = add_1472 + add_1483;
assign mul_1673 = slice_1667 * slice_1665;
assign slice_1862 = slice_1861[28:14];
assign slice_223 = mul_222[17:9];
assign concat_412 = {addW_410,slice_411};
assign add_601 = lsl_599 + mul_600;
assign slice_790 = slice_786[4:0];
assign slice_979 = slice_963[8:5];
assign slice_1168 = slice_1163[6:0];
assign slice_1357 = slice_1356[28:14];
assign mulnw_1546 = slice_1520 * slice_1545;
assign slice_1735 = addW_1719[17:0];
assign addW_1924 = slice_1864 + slice_1806;
assign slice_285 = mul_284[35:18];
assign add_474 = lsl_467 + add_473;
assign lsl_663 = add_662 << 5;
assign addW_852 = mul_850 + mul_851;
assign slice_1041 = addW_1025[8:0];
assign concat_1230 = {mul_1225,slice_1229};
assign slice_1419 = slice_1360[27:0];
assign mul_1608 = slice_1602 * slice_1600;
assign concat_1797 = {addW_1795,slice_1796};
assign mul_1986 = slice_1981 * slice_1952;
assign mulnw_158 = slice_157 * slice_123;
assign mul_347 = slice_343 * slice_346;
assign mulnw_536 = slice_510 * slice_496;
assign slice_725 = slice_721[6:0];
assign concat_914 = {addW_912,slice_913};
assign mul_1103 = slice_1101 * slice_1102;
assign mul_1292 = slice_1288 * slice_1291;
assign mul_1481 = slice_1476 * slice_1447;
assign slice_1670 = mul_1669[9:5];
assign slice_1859 = concat_1836[13:0];
assign slice_220 = addW_202[8:0];
assign addW_409 = add_397 + add_408;
assign add_598 = mulnw_596 + mulnw_597;
assign slice_787 = slice_786[9:5];
assign mul_976 = slice_952 * slice_972;
assign slice_1165 = slice_1148[13:0];
assign addW_1354 = slice_697 + slice_9;
assign lsl_1543 = mulnw_1542 << 10;
assign slice_1732 = mul_1725[5:0];
assign addW_1921 = slice_1861 + slice_1802;
assign slice_93 = slice_92[27:18];
assign slice_282 = slice_263[17:0];
assign lsl_471 = add_470 << 7;
assign slice_660 = slice_652[4:0];
assign concat_849 = {mul_844,slice_848};
assign slice_1038 = mul_1031[4:0];
assign slice_1227 = slice_1223[6:0];
assign slice_1416 = slice_1355[27:0];
assign slice_1605 = mul_1604[13:7];
assign subW_1794 = subW_1793 - concat_1713;
assign mulnw_1983 = slice_1978 * slice_1952;
assign mulnw_155 = slice_154 * slice_123;
assign slice_344 = slice_266[27:0];
assign mul_533 = slice_498 * slice_515;
assign slice_722 = slice_721[13:7];
assign subW_911 = subW_910 - mul_858;
assign mul_1100 = slice_1097 * slice_1099;
assign addW_1289 = slice_1282 + slice_1267;
assign mulnw_1478 = slice_1473 * slice_1447;
assign slice_1667 = slice_1661[4:0];
assign add_1856 = lsl_1849 + add_1855;
assign slice_28 = slice_16[6:0];
assign addW_217 = concat_213 + addW_216;
assign mul_406 = slice_401 * slice_372;
assign lsl_595 = mulnw_594 << 14;
assign slice_784 = slice_783[9:5];
assign mulnw_973 = slice_947 * slice_972;
assign concat_1162 = {addW_1160,slice_1161};
assign concat_1351 = {concat_696,slice_1350};
assign concat_1540 = {concat_1535,slice_1539};
assign mul_1729 = slice_1723 * slice_1721;
assign concat_1918 = {addW_1916,slice_1917};
assign addW_279 = concat_275 + addW_278;
assign mulnw_468 = slice_444 * slice_426;
assign mulnw_657 = slice_635 * slice_656;
assign slice_846 = slice_842[5:0];
assign mul_1035 = slice_1029 * slice_1027;
assign slice_1224 = slice_1223[13:7];
assign addW_1413 = concat_1393 + addW_1412;
assign slice_1602 = slice_1597[6:0];
assign slice_1791 = mul_1736[17:0];
assign lsl_1980 = mulnw_1979 << 10;
assign add_152 = lsl_150 + mul_151;
assign slice_341 = slice_262[27:0];
assign mulnw_530 = slice_492 * slice_515;
assign slice_719 = slice_699[13:0];
assign slice_908 = mul_881[8:0];
assign slice_1097 = slice_1096[13:7];
assign addW_1286 = slice_1281 + slice_1264;
assign lsl_1475 = mulnw_1474 << 10;
assign slice_1664 = addW_1663[18:9];
assign lsl_1853 = add_1852 << 7;
assign mul_25 = slice_18 * slice_24;
assign mul_214 = slice_204 * slice_210;
assign mulnw_403 = slice_398 * slice_372;
assign add_592 = lsl_590 + mul_591;
assign concat_781 = {concat_776,slice_780};
assign lsl_970 = mulnw_969 << 10;
assign addW_1159 = mul4_1157 + mul4_1158;
assign slice_1348 = concat_1140[55:0];
assign slice_1537 = addW_1521[8:0];
assign slice_1726 = mul_1725[11:6];
assign addW_1915 = add_1905 + add_1914;
assign slice_87 = slice_12[27:0];
assign mul_276 = slice_265 * slice_272;
assign add_465 = lsl_458 + add_464;
assign slice_654 = mul_653[17:9];
assign slice_843 = slice_842[11:6];
assign slice_1032 = mul_1031[9:5];
assign slice_1221 = slice_1203[13:0];
assign add_1410 = lsl_1408 + mul_1409;
assign slice_1599 = slice_1582[13:0];
assign subW_1788 = concat_1787 - concat_1733;
assign add_1977 = lsl_1969 + add_1976;
assign add_149 = mulnw_146 + mulnw_148;
assign addW_338 = concat_286 + subW_337;
assign mulnw_527 = slice_492 * slice_512;
assign addW_716 = concat_712 + addW_715;
assign add_905 = lsl_897 + add_904;
assign slice_1094 = mul_1087[6:0];
assign mul_1283 = slice_1281 * slice_1282;
assign add_1472 = lsl_1464 + add_1471;
assign slice_1661 = addW_1660[18:9];
assign mulnw_1850 = slice_1826 * slice_1808;
assign slice_22 = slice_21[56:28];
assign mul_211 = slice_209 * slice_210;
assign lsl_400 = mulnw_399 << 10;
assign add_589 = mulnw_587 + mulnw_588;
assign slice_778 = slice_762[17:0];
assign concat_967 = {concat_962,slice_966};
assign concat_1156 = {mul_1151,slice_1155};
assign subW_1345 = concat_1344 - concat_919;
assign slice_1534 = mul_1527[4:0];
assign slice_1723 = slice_1717[5:0];
assign mul_1912 = slice_1884 * slice_1869;
assign concat_84 = {addW_82,slice_83};
assign mul_273 = slice_271 * slice_272;
assign lsl_462 = add_461 << 7;
assign slice_651 = addW_633[8:0];
assign slice_840 = slice_839[11:6];
assign slice_1029 = slice_1023[4:0];
assign addW_1218 = concat_1214 + addW_1217;
assign add_1407 = mulnw_1405 + mulnw_1406;
assign concat_1596 = {addW_1594,slice_1595};
assign addW_1785 = concat_1761 + addW_1784;
assign lsl_1974 = add_1973 << 5;
assign mulnw_146 = slice_125 * slice_143;
assign concat_335 = {addW_333,slice_334};
assign concat_524 = {addW_522,slice_523};
assign mul4_713 = slice_701 * slice_709;
assign lsl_902 = add_901 << 5;
assign mul4_1091 = slice_1085 * slice_1083;
assign concat_1280 = {addW_1278,slice_1279};
assign lsl_1469 = add_1468 << 5;
assign slice_1658 = mul_1657[35:18];
assign add_1847 = lsl_1840 + add_1846;
assign mul_208 = slice_204 * slice_207;
assign add_397 = lsl_389 + add_396;
assign lsl_586 = mulnw_585 << 14;
assign slice_775 = mul_768[4:0];
assign slice_964 = addW_948[8:0];
assign slice_1153 = slice_1149[6:0];
assign addW_1342 = concat_1262 + subW_1341;
assign mul_1531 = slice_1525 * slice_1523;
assign slice_1720 = addW_1719[29:18];
assign mulnw_1909 = slice_1880 * slice_1869;
assign addW_81 = add_71 + add_80;
assign mul_270 = slice_265 * slice_269;
assign mulnw_459 = slice_428 * slice_442;
assign addW_648 = concat_644 + addW_647;
assign concat_837 = {concat_758,slice_836};
assign slice_1026 = addW_1025[18:9];
assign mul4_1215 = slice_1205 * slice_1211;
assign lsl_1404 = mulnw_1403 << 14;
assign addW_1593 = mul4_1591 + mul4_1592;
assign add_1782 = lsl_1780 + mul_1781;
assign slice_1971 = slice_1963[4:0];
assign slice_143 = slice_137[8:5];
assign addW_332 = add_320 + add_331;
assign addW_521 = mul_519 + mul_520;
assign mul_710 = slice_708 * slice_709;
assign mulnw_899 = slice_898 * slice_866;
assign slice_1088 = mul_1087[13:7];
assign addW_1277 = mul_1275 + mul_1276;
assign slice_1466 = slice_1458[4:0];
assign slice_1655 = slice_1637[17:0];
assign lsl_1844 = add_1843 << 7;
assign slice_16 = slice_14[28:14];
assign addW_205 = slice_198 + slice_183;
assign lsl_394 = add_393 << 5;
assign slice_583 = concat_582[27:14];
assign mul_772 = slice_766 * slice_764;
assign slice_961 = mul_954[4:0];
assign slice_1150 = slice_1149[14:7];
assign concat_1339 = {addW_1337,slice_1338};
assign slice_1528 = mul_1527[9:5];
assign slice_1717 = addW_1716[29:18];
assign mulnw_1906 = slice_1880 * slice_1866;
assign mul_78 = slice_47 * slice_29;
assign slice_267 = slice_266[55:28];
assign concat_456 = {concat_438,slice_455};
assign mul_645 = slice_635 * slice_641;
assign slice_834 = mul_779[17:0];
assign slice_1023 = addW_1022[18:9];
assign mul_1212 = slice_1210 * slice_1211;
assign add_1401 = lsl_1399 + mul_1400;
assign concat_1590 = {mul_1585,slice_1589};
assign add_1779 = mulnw_1777 + mulnw_1778;
assign mulnw_1968 = slice_1946 * slice_1967;
assign concat_140 = {concat_135,slice_139};
assign mul_329 = slice_324 * slice_295;
assign concat_518 = {mul_513,slice_517};
assign mul_707 = slice_701 * slice_706;
assign mulnw_896 = slice_895 * slice_866;
assign slice_1085 = slice_1079[6:0];
assign concat_1274 = {mul_1269,slice_1273};
assign mulnw_1463 = slice_1441 * slice_1462;
assign addW_1652 = concat_1648 + addW_1651;
assign mulnw_1841 = slice_1810 * slice_1824;
assign addW_202 = slice_197 + slice_180;
assign slice_391 = slice_383[4:0];
assign addW_580 = concat_576 + addW_579;
assign slice_769 = mul_768[9:5];
assign mul_958 = slice_952 * slice_950;
assign addW_1147 = slice_924 + slice_703;
assign subW_1336 = subW_1335 - mul_1283;
assign slice_1525 = slice_1519[4:0];
assign slice_1714 = concat_1713[55:28];
assign mul_1903 = slice_1868 * slice_1885;
assign mulnw_75 = slice_43 * slice_29;
assign slice_264 = slice_263[27:18];
assign slice_453 = mul_446[6:0];
assign mul_642 = slice_640 * slice_641;
assign subW_831 = concat_830 - concat_776;
assign slice_1020 = mul_1019[35:18];
assign mul_1209 = slice_1205 * slice_1208;
assign add_1398 = mulnw_1396 + mulnw_1397;
assign slice_1587 = slice_1583[6:0];
assign slice_1776 = slice_1757[4:0];
assign slice_1965 = mul_1964[17:9];
assign slice_137 = addW_121[8:0];
assign mulnw_326 = slice_321 * slice_295;
assign slice_515 = slice_511[6:0];
assign slice_704 = slice_703[56:28];
assign add_893 = lsl_891 + mul_892;
assign slice_1082 = addW_1081[28:14];
assign slice_1271 = slice_1267[5:0];
assign slice_1460 = mul_1459[17:9];
assign mul_1649 = slice_1639 * slice_1645;
assign concat_1838 = {concat_1820,slice_1837};
assign mul_199 = slice_197 * slice_198;
assign mulnw_388 = slice_366 * slice_387;
assign mul_577 = slice_568 * slice_573;
assign slice_766 = slice_760[4:0];
assign slice_955 = mul_954[9:5];
assign slice_1144 = addW_1143[57:29];
assign slice_1333 = mul_1306[8:0];
assign slice_1522 = addW_1521[18:9];
assign addW_1711 = concat_1659 + subW_1710;
assign mulnw_1900 = slice_1863 * slice_1885;
assign mulnw_72 = slice_43 * slice_24;
assign mul_450 = slice_444 * slice_442;
assign mul_639 = slice_635 * slice_638;
assign addW_828 = concat_804 + addW_827;
assign slice_1017 = slice_999[17:0];
assign slice_1206 = addW_1147[28:0];
assign lsl_1395 = mulnw_1394 << 14;
assign slice_1584 = slice_1583[14:7];
assign slice_1773 = slice_1757[8:5];
assign slice_1962 = addW_1944[8:0];
assign slice_134 = mul_127[4:0];
assign lsl_323 = mulnw_322 << 10;
assign slice_512 = slice_511[13:7];
assign slice_701 = slice_700[14:7];
assign add_890 = mulnw_887 + mulnw_889;
assign slice_1079 = addW_1078[28:14];
assign slice_1268 = slice_1267[11:6];
assign slice_1457 = addW_1439[8:0];
assign mul_1646 = slice_1644 * slice_1645;
assign slice_1835 = mul_1828[6:0];
assign concat_196 = {addW_194,slice_195};
assign slice_385 = mul_384[17:9];
assign mul_574 = slice_572 * slice_573;
assign slice_763 = slice_762[27:18];
assign slice_952 = slice_946[4:0];
assign slice_1141 = concat_1140[111:56];
assign add_1330 = lsl_1322 + add_1329;
assign slice_1519 = addW_1518[18:9];
assign concat_1708 = {addW_1706,slice_1707};
assign mulnw_1897 = slice_1863 * slice_1882;
assign mul_69 = slice_28 * slice_48;
assign addW_258 = concat_176 + subW_257;
assign slice_447 = mul_446[13:7];
assign addW_636 = slice_629 + slice_614;
assign add_825 = lsl_823 + mul_824;
assign addW_1014 = concat_1010 + addW_1013;
assign slice_1203 = addW_1143[28:0];
assign slice_1392 = concat_1391[27:14];
assign slice_1581 = addW_1359[56:0];
assign mul_1770 = slice_1746 * slice_1766;
assign addW_1959 = concat_1955 + addW_1958;
assign mul_131 = slice_125 * slice_123;
assign add_320 = lsl_312 + add_319;
assign slice_509 = slice_490[13:0];
assign slice_698 = slice_697[112:56];
assign mulnw_887 = slice_868 * slice_884;
assign slice_1076 = concat_1075[55:28];
assign slice_1265 = slice_1264[11:6];
assign addW_1454 = concat_1450 + addW_1453;
assign mul_1643 = slice_1639 * slice_1642;
assign mul_1832 = slice_1826 * slice_1824;
assign addW_193 = mul_191 + mul_192;
assign slice_382 = addW_364[8:0];
assign mul_571 = slice_568 * slice_570;
assign slice_760 = slice_759[27:18];
assign slice_949 = addW_948[18:9];
assign addW_1138 = concat_1077 + subW_1137;
assign lsl_1327 = add_1326 << 5;
assign slice_1516 = mul_1515[35:18];
assign addW_1705 = add_1693 + add_1704;
assign concat_1894 = {addW_1892,slice_1893};
assign mulnw_66 = slice_18 * slice_48;
assign concat_255 = {addW_253,slice_254};
assign slice_444 = slice_439[6:0];
assign addW_633 = slice_628 + slice_611;
assign add_822 = mulnw_820 + mulnw_821;
assign mul_1011 = slice_1001 * slice_1007;
assign addW_1200 = concat_1180 + addW_1199;
assign addW_1389 = concat_1385 + addW_1388;
assign slice_1578 = slice_1577[56:28];
assign mulnw_1767 = slice_1741 * slice_1766;
assign mul_1956 = slice_1946 * slice_1952;
assign slice_128 = mul_127[9:5];
assign lsl_317 = add_316 << 5;
assign addW_506 = concat_502 + addW_505;
assign slice_695 = concat_483[55:0];
assign slice_884 = slice_880[8:5];
assign addW_1073 = concat_1021 + subW_1072;
assign concat_1262 = {concat_1202,slice_1261};
assign mul_1451 = slice_1441 * slice_1447;
assign slice_1640 = slice_1581[27:0];
assign slice_1829 = mul_1828[13:7];
assign concat_190 = {mul_185,slice_189};
assign addW_379 = concat_375 + addW_378;
assign slice_568 = slice_567[13:7];
assign slice_757 = concat_734[13:0];
assign slice_946 = addW_945[18:9];
assign concat_1135 = {addW_1133,slice_1134};
assign mulnw_1324 = slice_1323 * slice_1291;
assign slice_1513 = addW_1495[17:0];
assign mul_1702 = slice_1697 * slice_1668;
assign addW_1891 = mul_1889 + mul_1890;
assign mulnw_63 = slice_18 * slice_45;
assign subW_252 = subW_251 - mul_199;
assign slice_441 = addW_424[13:0];
assign mul_630 = slice_628 * slice_629;
assign slice_819 = slice_800[4:0];
assign mul_1008 = slice_1006 * slice_1007;
assign add_1197 = lsl_1195 + mul_1196;
assign mul_1386 = slice_1377 * slice_1382;
assign slice_1575 = concat_1492[27:0];
assign lsl_1764 = mulnw_1763 << 10;
assign mul_1953 = slice_1951 * slice_1952;
assign slice_125 = slice_119[4:0];
assign slice_314 = slice_306[4:0];
assign mul4_503 = slice_492 * slice_499;
assign subW_692 = concat_691 - concat_260;
assign mul_881 = slice_879 * slice_880;
assign concat_1070 = {addW_1068,slice_1069};
assign slice_1259 = concat_1236[13:0];
assign mul_1448 = slice_1446 * slice_1447;
assign slice_1637 = slice_1577[27:0];
assign slice_1826 = slice_1821[6:0];
assign slice_187 = slice_183[5:0];
assign mul_376 = slice_366 * slice_372;
assign slice_565 = mul_558[6:0];
assign add_754 = lsl_747 + add_753;
assign slice_943 = mul_942[35:18];
assign addW_1132 = add_1122 + add_1131;
assign mulnw_1321 = slice_1320 * slice_1291;
assign addW_1510 = concat_1506 + addW_1509;
assign mulnw_1699 = slice_1694 * slice_1668;
assign concat_1888 = {mul_1883,slice_1887};
assign slice_60 = concat_58[27:14];
assign slice_249 = mul_222[8:0];
assign concat_438 = {addW_436,slice_437};
assign concat_627 = {addW_625,slice_626};
assign slice_816 = slice_800[8:5];
assign mul_1005 = slice_1001 * slice_1004;
assign add_1194 = mulnw_1192 + mulnw_1193;
assign mul_1383 = slice_1381 * slice_1382;
assign subW_1572 = concat_1571 - concat_1415;
assign concat_1761 = {concat_1756,slice_1760};
assign mul_1950 = slice_1946 * slice_1949;
assign slice_122 = addW_121[18:9];
assign mulnw_311 = slice_289 * slice_310;
assign mul_500 = slice_498 * slice_499;
assign addW_689 = concat_608 + subW_688;
assign concat_878 = {addW_876,slice_877};
assign addW_1067 = add_1055 + add_1066;
assign add_1256 = lsl_1249 + add_1255;
assign mul_1445 = slice_1441 * slice_1444;
assign addW_1634 = concat_1614 + addW_1633;
assign slice_1823 = slice_1806[13:0];
assign concat_2012 = {addW_2010,slice_2011};
assign slice_184 = slice_183[11:6];
assign mul_373 = slice_371 * slice_372;
assign mul4_562 = slice_556 * slice_554;
assign lsl_751 = add_750 << 7;
assign slice_940 = slice_921[17:0];
assign mul_1129 = slice_1101 * slice_1086;
assign add_1318 = lsl_1316 + mul_1317;
assign mul_1507 = slice_1497 * slice_1503;
assign lsl_1696 = mulnw_1695 << 10;
assign slice_1885 = slice_1881[6:0];
assign slice_57 = mul_49[6:0];
assign add_246 = lsl_238 + add_245;
assign addW_435 = mul4_433 + mul4_434;
assign addW_624 = mul_622 + mul_623;
assign mul_813 = slice_789 * slice_809;
assign slice_1002 = slice_924[27:0];
assign lsl_1191 = mulnw_1190 << 14;
assign mul_1380 = slice_1377 * slice_1379;
assign addW_1569 = concat_1517 + subW_1568;
assign slice_1758 = addW_1742[8:0];
assign addW_1947 = slice_1940 + slice_1925;
assign slice_119 = addW_118[18:9];
assign slice_308 = mul_307[17:9];
assign mul_497 = slice_492 * slice_496;
assign concat_686 = {addW_684,slice_685};
assign addW_875 = mul_873 + mul_874;
assign mul_1064 = slice_1059 * slice_1030;
assign lsl_1253 = add_1252 << 7;
assign addW_1442 = slice_1435 + slice_1420;
assign add_1631 = lsl_1629 + mul_1630;
assign concat_1820 = {addW_1818,slice_1819};
assign subW_2009 = subW_2008 - concat_1349;
assign slice_181 = slice_180[11:6];
assign mul_370 = slice_366 * slice_369;
assign slice_559 = mul_558[13:7];
assign mulnw_748 = slice_724 * slice_706;
assign addW_937 = concat_933 + addW_936;
assign mulnw_1126 = slice_1097 * slice_1086;
assign add_1315 = mulnw_1312 + mulnw_1314;
assign mul_1504 = slice_1502 * slice_1503;
assign add_1693 = lsl_1685 + add_1692;
assign slice_1882 = slice_1881[13:7];
assign mul_54 = slice_47 * slice_45;
assign lsl_243 = add_242 << 5;
assign concat_432 = {mul_427,slice_431};
assign concat_621 = {mul_616,slice_620};
assign mulnw_810 = slice_784 * slice_809;
assign slice_999 = slice_920[27:0];
assign add_1188 = lsl_1186 + mul_1187;
assign slice_1377 = slice_1376[13:7];
assign concat_1566 = {addW_1564,slice_1565};
assign slice_1755 = mul_1748[4:0];
assign addW_1944 = slice_1939 + slice_1922;
assign slice_305 = addW_287[8:0];
assign slice_494 = addW_493[57:29];
assign subW_683 = subW_682 - mul_630;
assign concat_872 = {mul_867,slice_871};
assign mulnw_1061 = slice_1056 * slice_1030;
assign mulnw_1250 = slice_1226 * slice_1208;
assign addW_1439 = slice_1434 + slice_1417;
assign add_1628 = mulnw_1626 + mulnw_1627;
assign addW_1817 = mul4_1815 + mul4_1816;
assign slice_2006 = concat_1797[56:0];
assign addW_367 = slice_360 + slice_345;
assign slice_556 = slice_550[6:0];
assign add_745 = lsl_738 + add_744;
assign mul_934 = slice_923 * slice_930;
assign mulnw_1123 = slice_1097 * slice_1083;
assign mulnw_1312 = slice_1293 * slice_1309;
assign mul_1501 = slice_1497 * slice_1500;
assign lsl_1690 = add_1689 << 5;
assign slice_1879 = slice_1861[13:0];
assign concat_51 = {mul_46,slice_50};
assign mulnw_240 = slice_239 * slice_207;
assign slice_429 = slice_425[6:0];
assign slice_618 = slice_614[5:0];
assign lsl_807 = mulnw_806 << 10;
assign addW_996 = concat_944 + subW_995;
assign add_1185 = mulnw_1183 + mulnw_1184;
assign slice_1374 = mul_1367[6:0];
assign addW_1563 = add_1551 + add_1562;
assign mul_1752 = slice_1746 * slice_1744;
assign mul_1941 = slice_1939 * slice_1940;
assign addW_302 = concat_298 + addW_301;
assign slice_491 = slice_490[28:14];
assign slice_680 = mul_653[8:0];
assign slice_869 = slice_865[4:0];
assign lsl_1058 = mulnw_1057 << 10;
assign add_1247 = lsl_1240 + add_1246;
assign mul_1436 = slice_1434 * slice_1435;
assign lsl_1625 = mulnw_1624 << 14;
assign concat_1814 = {mul_1809,slice_1813};
assign subW_2003 = concat_2002 - concat_1576;
assign slice_175 = concat_173[55:28];
assign addW_364 = slice_359 + slice_342;
assign slice_553 = slice_552[28:14];
assign lsl_742 = add_741 << 7;
assign mul_931 = slice_929 * slice_930;
assign mul_1120 = slice_1085 * slice_1102;
assign slice_1309 = slice_1305[8:5];
assign addW_1498 = slice_1419 + slice_1361;
assign slice_1687 = slice_1679[4:0];
assign addW_1876 = concat_1872 + addW_1875;
assign slice_48 = slice_44[6:0];
assign mulnw_237 = slice_236 * slice_207;
assign slice_426 = slice_425[14:7];
assign slice_615 = slice_614[11:6];
assign concat_804 = {concat_799,slice_803};
assign concat_993 = {addW_991,slice_992};
assign lsl_1182 = mulnw_1181 << 14;
assign mul4_1371 = slice_1365 * slice_1363;
assign mul_1560 = slice_1555 * slice_1526;
assign slice_1749 = mul_1748[9:5];
assign concat_1938 = {addW_1936,slice_1937};
assign slice_110 = slice_87[17:0];
assign mul_299 = slice_289 * slice_295;
assign add_677 = lsl_669 + add_676;
assign slice_866 = slice_865[9:5];
assign add_1055 = lsl_1047 + add_1054;
assign lsl_1244 = add_1243 << 7;
assign concat_1433 = {addW_1431,slice_1432};
assign add_1622 = lsl_1620 + mul_1621;
assign slice_1811 = slice_1807[6:0];
assign addW_2000 = concat_1920 + subW_1999;
assign slice_172 = mul_112[17:0];
assign mul_361 = slice_359 * slice_360;
assign slice_550 = slice_549[28:14];
assign mulnw_739 = slice_708 * slice_722;
assign mul_928 = slice_923 * slice_927;
assign mulnw_1117 = slice_1080 * slice_1102;
assign mul_1306 = slice_1304 * slice_1305;
assign addW_1495 = slice_1416 + slice_1356;
assign mulnw_1684 = slice_1662 * slice_1683;
assign mul4_1873 = slice_1863 * slice_1869;
assign slice_45 = slice_44[13:7];
assign add_234 = lsl_232 + mul_233;
assign slice_423 = slice_422[14:7];
assign slice_612 = slice_611[11:6];
assign slice_801 = addW_785[8:0];
assign addW_990 = add_978 + add_989;
assign slice_1179 = concat_1178[27:14];
assign slice_1368 = mul_1367[13:7];
assign mulnw_1557 = slice_1552 * slice_1526;
assign slice_1746 = slice_1740[4:0];
assign addW_1935 = mul_1933 + mul_1934;
assign slice_107 = mul_99[4:0];
assign mul_296 = slice_294 * slice_295;
assign slice_485 = concat_483[111:56];
assign lsl_674 = add_673 << 5;
assign slice_863 = slice_862[9:5];
assign lsl_1052 = add_1051 << 5;
assign mulnw_1241 = slice_1210 * slice_1224;
assign addW_1430 = mul_1428 + mul_1429;
assign add_1619 = mulnw_1617 + mulnw_1618;
assign slice_1808 = slice_1807[14:7];
assign concat_1997 = {addW_1995,slice_1996};
assign subW_169 = concat_168 - concat_108;
assign concat_358 = {addW_356,slice_357};
assign slice_547 = concat_524[13:0];
assign concat_736 = {concat_718,slice_735};
assign slice_925 = slice_924[55:28];
assign mulnw_1114 = slice_1080 * slice_1099;
assign concat_1303 = {addW_1301,slice_1302};
assign concat_1492 = {addW_1490,slice_1491};
assign slice_1681 = mul_1680[17:9];
assign mul_1870 = slice_1868 * slice_1869;
assign slice_42 = slice_14[13:0];
assign add_231 = mulnw_228 + mulnw_230;
assign slice_798 = mul_791[4:0];
assign mul_987 = slice_982 * slice_953;
assign addW_1176 = concat_1172 + addW_1175;
assign slice_1365 = slice_1357[6:0];
assign lsl_1554 = mulnw_1553 << 10;
assign slice_1743 = addW_1742[18:9];
assign concat_1932 = {mul_1927,slice_1931};
assign mul_104 = slice_97 * slice_94;
assign mul_293 = slice_289 * slice_292;
assign slice_482 = concat_417[27:0];
assign mulnw_671 = slice_670 * slice_638;
assign concat_860 = {concat_855,slice_859};
assign slice_1049 = slice_1041[4:0];
assign concat_1238 = {concat_1220,slice_1237};
assign concat_1427 = {mul_1422,slice_1426};
assign lsl_1616 = mulnw_1615 << 14;
assign addW_1805 = slice_1581 + slice_1360;
assign subW_1994 = subW_1993 - mul_1941;
assign addW_166 = concat_140 + addW_165;
assign addW_355 = mul_353 + mul_354;
assign add_544 = lsl_537 + add_543;
assign slice_733 = mul_726[6:0];
assign slice_922 = slice_921[27:18];
assign concat_1111 = {addW_1109,slice_1110};
assign addW_1300 = mul_1298 + mul_1299;
assign subW_1489 = subW_1488 - mul_1436;
assign slice_1678 = addW_1660[8:0];
assign mul_1867 = slice_1863 * slice_1866;
assign slice_39 = mul_30[6:0];
assign mulnw_228 = slice_209 * slice_225;
assign concat_417 = {addW_415,slice_416};
assign concat_606 = {addW_604,slice_605};
assign mul_795 = slice_789 * slice_787;
assign mulnw_984 = slice_979 * slice_953;
assign mul_1173 = slice_1164 * slice_1169;
assign slice_1362 = slice_1361[28:14];
assign add_1551 = lsl_1543 + add_1550;
assign slice_1740 = addW_1739[18:9];
assign slice_1929 = slice_1925[5:0];
assign concat_101 = {mul_95,slice_100};
assign addW_290 = slice_283 + slice_268;
assign subW_479 = concat_478 - concat_340;
assign mulnw_668 = slice_667 * slice_638;
assign slice_857 = addW_841[17:0];
assign mulnw_1046 = slice_1024 * slice_1045;
assign slice_1235 = mul_1228[6:0];
assign slice_1424 = slice_1420[4:0];
assign slice_1613 = concat_1612[27:14];
assign slice_1802 = addW_1801[57:29];
assign slice_1991 = mul_1964[8:0];
assign add_163 = lsl_161 + mul_162;
assign concat_352 = {mul_347,slice_351};
assign lsl_541 = add_540 << 7;
assign mul_730 = slice_724 * slice_722;
assign concat_919 = {addW_917,slice_918};
assign addW_1108 = mul_1106 + mul_1107;
assign concat_1297 = {mul_1292,slice_1296};
assign slice_1486 = mul_1459[8:0];
assign addW_1675 = concat_1671 + addW_1674;
assign slice_1864 = addW_1805[28:0];
assign mul4_36 = slice_28 * slice_24;
assign slice_225 = slice_221[8:5];
assign subW_414 = subW_413 - mul_361;
assign addW_603 = add_593 + add_602;
assign slice_792 = mul_791[9:5];
assign lsl_981 = mulnw_980 << 10;
assign mul_1170 = slice_1168 * slice_1169;
assign addW_1359 = slice_702 + slice_20;
assign lsl_1548 = add_1547 << 5;
assign slice_1737 = mul_1736[35:18];
assign slice_1926 = slice_1925[11:6];
assign slice_98 = slice_93[4:0];
assign addW_287 = slice_282 + slice_264;
assign addW_476 = concat_456 + addW_475;
assign add_665 = lsl_663 + mul_664;
assign slice_854 = mul_847[5:0];
assign slice_1043 = mul_1042[17:9];
assign mul_1232 = slice_1226 * slice_1224;
assign slice_1421 = slice_1420[9:5];
assign addW_1610 = concat_1606 + addW_1609;
assign concat_1799 = {concat_1576,slice_1798};
assign add_1988 = lsl_1980 + add_1987;
assign add_160 = mulnw_158 + mulnw_159;
assign slice_349 = slice_345[4:0];
assign mulnw_538 = slice_514 * slice_496;
assign slice_727 = mul_726[13:7];
assign subW_916 = subW_915 - concat_835;
assign concat_1105 = {mul_1100,slice_1104};
assign slice_1294 = slice_1290[4:0];
assign add_1483 = lsl_1475 + add_1482;
assign mul_1672 = slice_1662 * slice_1668;
assign slice_1861 = addW_1801[28:0];
assign concat_33 = {mul_25,slice_32};
assign mul_222 = slice_220 * slice_221;
assign slice_411 = mul_384[8:0];
assign mul_600 = slice_572 * slice_557;
assign slice_789 = slice_783[4:0];
assign add_978 = lsl_970 + add_977;
assign mul_1167 = slice_1164 * slice_1166;
assign slice_1356 = slice_1355[56:28];
assign slice_1545 = slice_1537[4:0];
assign slice_1734 = addW_1716[17:0];
assign slice_1923 = slice_1922[11:6];
assign mul_95 = slice_91 * slice_94;
assign mul_284 = slice_282 * slice_283;
assign add_473 = lsl_471 + mul_472;
assign add_662 = mulnw_659 + mulnw_661;
assign mul_851 = slice_845 * slice_843;
assign slice_1040 = addW_1022[8:0];
assign slice_1229 = mul_1228[13:7];
assign slice_1418 = slice_1417[9:5];
assign mul_1607 = slice_1598 * slice_1603;
assign slice_1796 = concat_1713[27:0];
assign lsl_1985 = add_1984 << 5;
assign slice_157 = slice_136[4:0];
assign slice_346 = slice_345[9:5];
assign add_535 = lsl_528 + add_534;
assign slice_724 = slice_719[6:0];
assign slice_913 = mul_858[17:0];
assign slice_1102 = slice_1098[6:0];
assign slice_1291 = slice_1290[9:5];
assign lsl_1480 = add_1479 << 5;
assign mul_1669 = slice_1667 * slice_1668;
assign addW_1858 = concat_1838 + addW_1857;
assign mul_30 = slice_28 * slice_29;
assign concat_219 = {addW_217,slice_218};
assign add_408 = lsl_400 + add_407;
assign mulnw_597 = slice_568 * slice_557;
assign slice_786 = addW_785[18:9];
assign lsl_975 = add_974 << 5;
assign slice_1164 = slice_1163[13:7];
assign mulnw_1542 = slice_1520 * slice_1541;
assign addW_1731 = concat_1727 + addW_1730;
assign concat_1920 = {concat_1860,slice_1919};
assign slice_92 = slice_21[27:0];
assign concat_281 = {addW_279,slice_280};
assign add_470 = mulnw_468 + mulnw_469;
assign mulnw_659 = slice_640 * slice_656;
assign slice_848 = mul_847[11:6];
assign addW_1037 = concat_1033 + addW_1036;
assign slice_1226 = slice_1221[6:0];
assign concat_1415 = {addW_1413,slice_1414};
assign mul_1604 = slice_1602 * slice_1603;
assign subW_1793 = concat_1792 - concat_1636;
assign mulnw_1982 = slice_1981 * slice_1949;
assign slice_154 = slice_136[8:5];
assign slice_343 = slice_342[9:5];
assign lsl_532 = add_531 << 7;
assign slice_721 = slice_704[13:0];
assign subW_910 = concat_909 - concat_855;
assign slice_1099 = slice_1098[13:7];
assign slice_1288 = slice_1287[9:5];
assign mulnw_1477 = slice_1476 * slice_1444;
assign mul_1666 = slice_1662 * slice_1665;
assign add_1855 = lsl_1853 + mul_1854;
assign addW_216 = mul_214 + mul_215;
assign lsl_405 = add_404 << 5;
assign mulnw_594 = slice_568 * slice_554;
assign slice_783 = addW_782[18:9];
assign slice_972 = slice_964[4:0];
assign slice_1161 = mul_1154[6:0];
assign slice_1350 = concat_1349[225:113];
assign slice_1539 = mul_1538[17:9];
assign mul_1728 = slice_1718 * slice_1724;
assign slice_1917 = concat_1894[13:0];
assign slice_89 = slice_87[27:18];
assign addW_278 = mul_276 + mul_277;
assign lsl_467 = mulnw_466 << 14;
assign slice_656 = slice_652[8:5];
assign slice_845 = slice_839[5:0];
assign mul_1034 = slice_1024 * slice_1030;
assign slice_1223 = slice_1206[13:0];
assign addW_1412 = add_1402 + add_1411;
assign mul_1601 = slice_1598 * slice_1600;
assign addW_1790 = concat_1738 + subW_1789;
assign mulnw_1979 = slice_1978 * slice_1949;
assign mul_151 = slice_125 * slice_147;
assign concat_340 = {addW_338,slice_339};
assign mulnw_529 = slice_498 * slice_512;
assign concat_718 = {addW_716,slice_717};
assign addW_907 = concat_883 + addW_906;
assign slice_1096 = addW_1078[13:0];
assign concat_1285 = {concat_1280,slice_1284};
assign mulnw_1474 = slice_1473 * slice_1444;
assign addW_1663 = slice_1656 + slice_1641;
assign add_1852 = mulnw_1850 + mulnw_1851;
assign slice_24 = slice_23[14:7];
assign concat_213 = {mul_208,slice_212};
assign mulnw_402 = slice_401 * slice_369;
assign mul_591 = slice_556 * slice_573;
assign slice_780 = mul_779[35:18];
assign mulnw_969 = slice_947 * slice_968;
assign mul4_1158 = slice_1152 * slice_1150;
assign addW_1347 = concat_1142 + subW_1346;
assign slice_1536 = addW_1518[8:0];
assign mul_1725 = slice_1723 * slice_1724;
assign add_1914 = lsl_1907 + add_1913;
assign concat_275 = {mul_270,slice_274};
assign add_464 = lsl_462 + mul_463;
assign mul_653 = slice_651 * slice_652;
assign slice_842 = addW_841[29:18];
assign mul_1031 = slice_1029 * slice_1030;
assign concat_1220 = {addW_1218,slice_1219};
assign mul_1409 = slice_1381 * slice_1366;
assign slice_1598 = slice_1597[13:7];
assign concat_1787 = {addW_1785,slice_1786};
assign add_1976 = lsl_1974 + mul_1975;
assign mulnw_148 = slice_120 * slice_147;
assign subW_337 = subW_336 - mul_284;
assign concat_526 = {concat_508,slice_525};
assign addW_715 = mul4_713 + mul4_714;
assign add_904 = lsl_902 + mul_903;
assign addW_1093 = concat_1089 + addW_1092;
assign slice_1282 = addW_1266[17:0];
assign add_1471 = lsl_1469 + mul_1470;
assign addW_1660 = slice_1655 + slice_1638;
assign lsl_1849 = mulnw_1848 << 14;
assign slice_21 = slice_20[112:56];
assign slice_210 = slice_206[4:0];
assign mulnw_399 = slice_398 * slice_369;
assign mulnw_588 = slice_551 * slice_573;
assign slice_777 = slice_759[17:0];
assign slice_966 = mul_965[17:9];
assign slice_1155 = mul_1154[13:7];
assign concat_1344 = {addW_1342,slice_1343};
assign addW_1533 = concat_1529 + addW_1532;
assign mul_1722 = slice_1718 * slice_1721;
assign lsl_1911 = add_1910 << 7;
assign slice_83 = concat_58[13:0];
assign slice_272 = slice_268[4:0];
assign add_461 = mulnw_459 + mulnw_460;
assign concat_650 = {addW_648,slice_649};
assign slice_839 = addW_838[29:18];
assign mul_1028 = slice_1024 * slice_1027;
assign addW_1217 = mul4_1215 + mul4_1216;
assign mulnw_1406 = slice_1377 * slice_1366;
assign slice_1595 = mul_1588[6:0];
assign addW_1784 = add_1772 + add_1783;
assign add_1973 = mulnw_1970 + mulnw_1972;
assign lsl_145 = mulnw_144 << 10;
assign slice_334 = mul_307[8:0];
assign slice_523 = mul_516[6:0];
assign concat_712 = {mul_707,slice_711};
assign add_901 = mulnw_899 + mulnw_900;
assign mul4_1090 = slice_1080 * slice_1086;
assign slice_1279 = mul_1272[5:0];
assign add_1468 = mulnw_1465 + mulnw_1467;
assign mul_1657 = slice_1655 * slice_1656;
assign add_1846 = lsl_1844 + mul_1845;
assign slice_18 = slice_16[14:7];
assign slice_207 = slice_206[9:5];
assign add_396 = lsl_394 + mul_395;
assign mulnw_585 = slice_551 * slice_570;
assign addW_774 = concat_770 + addW_773;
assign slice_963 = addW_945[8:0];
assign slice_1152 = slice_1145[6:0];
assign subW_1341 = subW_1340 - concat_1260;
assign mul_1530 = slice_1520 * slice_1526;
assign addW_1719 = slice_1640 + slice_1582;
assign mulnw_1908 = slice_1884 * slice_1866;
assign add_80 = lsl_73 + add_79;
assign slice_269 = slice_268[9:5];
assign lsl_458 = mulnw_457 << 14;
assign addW_647 = mul_645 + mul_646;
assign slice_836 = concat_835[55:28];
assign addW_1025 = slice_1018 + slice_1003;
assign concat_1214 = {mul_1209,slice_1213};
assign mulnw_1403 = slice_1377 * slice_1363;
assign mul4_1592 = slice_1586 * slice_1584;
assign mul_1781 = slice_1776 * slice_1747;
assign mulnw_1970 = slice_1951 * slice_1967;
assign add_331 = lsl_323 + add_330;
assign mul_520 = slice_514 * slice_512;
assign slice_709 = slice_705[6:0];
assign slice_898 = slice_879[4:0];
assign mul_1087 = slice_1085 * slice_1086;
assign mul_1276 = slice_1270 * slice_1268;
assign mulnw_1465 = slice_1446 * slice_1462;
assign concat_1654 = {addW_1652,slice_1653};
assign add_1843 = mulnw_1841 + mulnw_1842;
assign slice_204 = slice_203[9:5];
assign add_393 = mulnw_390 + mulnw_392;
assign concat_582 = {addW_580,slice_581};
assign mul_771 = slice_761 * slice_767;
assign addW_960 = concat_956 + addW_959;
assign slice_1149 = slice_1148[28:14];
assign slice_1338 = mul_1283[17:0];
assign mul_1527 = slice_1525 * slice_1526;
assign addW_1716 = slice_1637 + slice_1578;
assign add_1905 = lsl_1898 + add_1904;
assign lsl_77 = add_76 << 7;
assign slice_266 = slice_20[55:0];
assign slice_455 = concat_454[27:14];
assign concat_644 = {mul_639,slice_643};
assign addW_833 = concat_781 + subW_832;
assign addW_1022 = slice_1017 + slice_1000;
assign slice_1211 = slice_1207[6:0];
assign mul_1400 = slice_1365 * slice_1382;
assign slice_1589 = mul_1588[13:7];
assign mulnw_1778 = slice_1773 * slice_1747;
assign slice_1967 = slice_1963[8:5];
assign slice_139 = mul_138[17:9];
assign lsl_328 = add_327 << 5;
assign slice_517 = mul_516[13:7];
assign slice_706 = slice_705[14:7];
assign slice_895 = slice_879[8:5];
assign mul_1084 = slice_1080 * slice_1083;
assign slice_1273 = mul_1272[11:6];
assign slice_1462 = slice_1458[8:5];
assign addW_1651 = mul_1649 + mul_1650;
assign lsl_1840 = mulnw_1839 << 14;
assign slice_12 = slice_9[112:56];
assign concat_201 = {concat_196,slice_200};
assign mulnw_390 = slice_371 * slice_387;
assign addW_579 = mul_577 + mul_578;
assign mul_768 = slice_766 * slice_767;
assign mul_957 = slice_947 * slice_953;
assign slice_1146 = slice_1145[14:7];
assign subW_1335 = concat_1334 - concat_1280;
assign mul_1524 = slice_1520 * slice_1523;
assign concat_1713 = {addW_1711,slice_1712};
assign lsl_1902 = add_1901 << 7;
assign mulnw_74 = slice_47 * slice_24;
assign slice_263 = slice_262[55:28];
assign addW_452 = concat_448 + addW_451;
assign slice_641 = slice_637[4:0];
assign concat_830 = {addW_828,slice_829};
assign mul_1019 = slice_1017 * slice_1018;
assign slice_1208 = slice_1207[14:7];
assign mulnw_1397 = slice_1358 * slice_1382;
assign slice_1586 = slice_1579[6:0];
assign lsl_1775 = mulnw_1774 << 10;
assign mul_1964 = slice_1962 * slice_1963;
assign slice_136 = addW_118[8:0];
assign mulnw_325 = slice_324 * slice_292;
assign slice_514 = slice_509[6:0];
assign slice_703 = slice_702[112:56];
assign mul_892 = slice_868 * slice_888;
assign addW_1081 = slice_1002 + slice_925;
assign slice_1270 = slice_1264[5:0];
assign mul_1459 = slice_1457 * slice_1458;
assign concat_1648 = {mul_1643,slice_1647};
assign slice_1837 = concat_1836[27:14];
assign slice_9 = IN1[225:113];
assign slice_198 = addW_182[17:0];
assign slice_387 = slice_383[8:5];
assign concat_576 = {mul_571,slice_575};
assign mul_765 = slice_761 * slice_764;
assign mul_954 = slice_952 * slice_953;
assign addW_1143 = slice_920 + slice_698;
assign addW_1332 = concat_1308 + addW_1331;
assign addW_1521 = slice_1514 + slice_1499;
assign subW_1710 = subW_1709 - mul_1657;
assign mulnw_1899 = slice_1868 * slice_1882;
assign add_71 = lsl_64 + add_70;
assign concat_260 = {addW_258,slice_259};
assign mul_449 = slice_440 * slice_445;
assign slice_638 = slice_637[9:5];
assign addW_827 = add_815 + add_826;
assign concat_1016 = {addW_1014,slice_1015};
assign slice_1205 = slice_1204[14:7];
assign mulnw_1394 = slice_1358 * slice_1379;
assign slice_1583 = slice_1582[28:14];
assign add_1772 = lsl_1764 + add_1771;
assign concat_1961 = {addW_1959,slice_1960};
assign addW_133 = concat_129 + addW_132;
assign mulnw_322 = slice_321 * slice_292;
assign slice_511 = slice_494[13:0];
assign slice_700 = slice_699[28:14];
assign mulnw_889 = slice_863 * slice_888;
assign addW_1078 = slice_999 + slice_921;
assign slice_1267 = addW_1266[29:18];
assign concat_1456 = {addW_1454,slice_1455};
assign slice_1645 = slice_1641[4:0];
assign addW_1834 = concat_1830 + addW_1833;
assign slice_195 = mul_188[5:0];
assign mul_384 = slice_382 * slice_383;
assign slice_573 = slice_569[6:0];
assign slice_762 = slice_703[27:0];
assign mul_951 = slice_947 * slice_950;
assign concat_1140 = {addW_1138,slice_1139};
assign add_1329 = lsl_1327 + mul_1328;
assign addW_1518 = slice_1513 + slice_1496;
assign slice_1707 = mul_1680[8:0];
assign concat_1896 = {concat_1878,slice_1895};
assign lsl_68 = add_67 << 7;
assign subW_257 = subW_256 - concat_173;
assign mul_446 = slice_444 * slice_445;
assign slice_635 = slice_634[9:5];
assign mul_824 = slice_819 * slice_790;
assign addW_1013 = mul_1011 + mul_1012;
assign concat_1202 = {addW_1200,slice_1201};
assign concat_1391 = {addW_1389,slice_1390};
assign slice_1580 = slice_1579[14:7];
assign lsl_1769 = add_1768 << 5;
assign addW_1958 = mul_1956 + mul_1957;
assign mul_130 = slice_120 * slice_126;
assign add_319 = lsl_317 + mul_318;
assign concat_508 = {addW_506,slice_507};
assign slice_697 = IN1[112:0];
assign lsl_886 = mulnw_885 << 10;
assign concat_1075 = {addW_1073,slice_1074};
assign slice_1264 = addW_1263[29:18];
assign addW_1453 = mul_1451 + mul_1452;
assign slice_1642 = slice_1641[9:5];
assign mul_1831 = slice_1822 * slice_1827;
assign mul_192 = slice_186 * slice_184;
assign concat_381 = {addW_379,slice_380};
assign slice_570 = slice_569[13:7];
assign slice_759 = slice_698[27:0];
assign addW_948 = slice_941 + slice_926;
assign subW_1137 = subW_1136 - concat_1075;
assign add_1326 = mulnw_1324 + mulnw_1325;
assign mul_1515 = slice_1513 * slice_1514;
assign add_1704 = lsl_1696 + add_1703;
assign slice_1893 = mul_1886[6:0];
assign mulnw_65 = slice_28 * slice_45;
assign slice_254 = mul_199[17:0];
assign mul_443 = slice_440 * slice_442;
assign concat_632 = {concat_627,slice_631};
assign mulnw_821 = slice_816 * slice_790;
assign concat_1010 = {mul_1005,slice_1009};
assign addW_1199 = add_1189 + add_1198;
assign addW_1388 = mul_1386 + mul_1387;
assign slice_1577 = addW_1354[56:0];
assign slice_1766 = slice_1758[4:0];
assign concat_1955 = {mul_1950,slice_1954};
assign mul_127 = slice_125 * slice_126;
assign add_316 = mulnw_313 + mulnw_315;
assign addW_505 = mul4_503 + mul4_504;
assign addW_694 = concat_486 + subW_693;
assign concat_883 = {concat_878,slice_882};
assign subW_1072 = subW_1071 - mul_1019;
assign slice_1261 = concat_1260[57:29];
assign concat_1450 = {mul_1445,slice_1449};
assign slice_1639 = slice_1638[9:5];
assign mul_1828 = slice_1826 * slice_1827;
assign OUTPUT = concat_2012;
    endmodule