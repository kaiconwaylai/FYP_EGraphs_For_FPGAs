//Alpha = 0.005. Cost: LUTs = 187110. DSPs = 0.  

`timescale 1ns / 1ps
    module mult(
        input[1023:0] IN1,
        input[1023:0] IN2,
        output[2047:0] OUTPUT
    );
wire [65:0] addW_4663;
wire [33:0] mul_756;
wire [33:0] add_5419;
wire [17:0] slice_1512;
wire [17:0] slice_6175;
wire [32:0] lsl_2268;
wire [7:0] slice_6931;
wire [25:0] lsl_3024;
wire [7:0] slice_3780;
wire [15:0] slice_4536;
wire [19:0] addW_629;
wire [15:0] mul_5292;
wire [51:0] addW_1385;
wire [15:0] mul_6048;
wire [17:0] add_2141;
wire [39:0] mul_6804;
wire [66:0] concat_2897;
wire [99:0] concat_7560;
wire [19:0] addW_3653;
wire [15:0] mul_4409;
wire [15:0] mul_502;
wire [31:0] slice_5165;
wire [65:0] concat_1258;
wire [17:0] slice_5921;
wire [45:0] concat_2014;
wire [15:0] mulnw_6677;
wire [31:0] slice_2770;
wire [13:0] slice_7433;
wire [8:0] slice_3526;
wire [70:0] subW_4282;
wire [7:0] slice_375;
wire [263:0] subW_5038;
wire [195:0] addW_1131;
wire [8:0] slice_5794;
wire [7:0] slice_1887;
wire [39:0] mul_6550;
wire [31:0] slice_2643;
wire [16:0] slice_7306;
wire [31:0] slice_3399;
wire [26:0] add_4155;
wire [25:0] lsl_248;
wire [19:0] addW_4911;
wire [31:0] mul_1004;
wire [47:0] addW_5667;
wire [98:0] concat_1760;
wire [131:0] concat_6423;
wire [17:0] slice_2516;
wire [15:0] slice_7179;
wire [7:0] slice_3272;
wire [17:0] slice_4028;
wire [68:0] subW_121;
wire [16:0] mulnw_4784;
wire [13:0] slice_877;
wire [33:0] add_5540;
wire [16:0] mulnw_1633;
wire [33:0] mul_6296;
wire [45:0] concat_2389;
wire [26:0] add_7052;
wire [98:0] concat_3145;
wire [63:0] slice_3901;
wire [130:0] concat_4657;
wire [66:0] addW_750;
wire [7:0] slice_5413;
wire [65:0] concat_1506;
wire [127:0] slice_6169;
wire [31:0] mul_2262;
wire [26:0] add_6925;
wire [32:0] lsl_3018;
wire [15:0] slice_3774;
wire [33:0] addW_4530;
wire [17:0] slice_623;
wire [7:0] slice_5286;
wire [49:0] concat_1379;
wire [7:0] slice_6042;
wire [16:0] mulnw_2135;
wire [17:0] slice_6798;
wire [15:0] mul_2891;
wire [33:0] add_7554;
wire [27:0] mul_3647;
wire [7:0] slice_4403;
wire [7:0] slice_496;
wire [41:0] subW_5159;
wire [19:0] addW_1252;
wire [19:0] addW_5915;
wire [13:0] slice_2008;
wire [8:0] slice_6671;
wire [34:0] addW_2764;
wire [33:0] add_7427;
wire [17:0] add_3520;
wire [39:0] mul_4276;
wire [26:0] add_369;
wire [133:0] concat_5032;
wire [71:0] subW_1125;
wire [33:0] mul_5788;
wire [15:0] slice_1881;
wire [17:0] slice_6544;
wire [31:0] slice_2637;
wire [128:0] slice_7300;
wire [41:0] subW_3393;
wire [16:0] mulnw_4149;
wire [32:0] lsl_242;
wire [31:0] mul_4905;
wire [16:0] slice_998;
wire [45:0] concat_5661;
wire [40:0] subW_1754;
wire [17:0] slice_6417;
wire [34:0] addW_2510;
wire [25:0] lsl_7173;
wire [15:0] slice_3266;
wire [19:0] addW_4022;
wire [33:0] add_115;
wire [33:0] add_4778;
wire [31:0] slice_871;
wire [7:0] slice_5534;
wire [7:0] slice_1627;
wire [31:0] slice_6290;
wire [13:0] slice_2383;
wire [16:0] mulnw_7046;
wire [40:0] subW_3139;
wire [99:0] addW_3895;
wire [15:0] slice_4651;
wire [31:0] slice_744;
wire [7:0] slice_5407;
wire [19:0] addW_1500;
wire [63:0] slice_6163;
wire [64:0] slice_2256;
wire [15:0] mulnw_6919;
wire [15:0] mul_3012;
wire [33:0] addW_3768;
wire [17:0] slice_4524;
wire [66:0] concat_617;
wire [15:0] slice_5280;
wire [15:0] slice_1373;
wire [15:0] slice_6036;
wire [25:0] lsl_2129;
wire [34:0] addW_6792;
wire [7:0] slice_2885;
wire [7:0] slice_7548;
wire [31:0] slice_3641;
wire [26:0] add_4397;
wire [15:0] slice_490;
wire [17:0] slice_5153;
wire [17:0] slice_1246;
wire [27:0] mul_5909;
wire [47:0] addW_2002;
wire [17:0] add_6665;
wire [15:0] mulnw_2758;
wire [7:0] slice_7421;
wire [16:0] mulnw_3514;
wire [17:0] slice_4270;
wire [15:0] mulnw_363;
wire [17:0] slice_5026;
wire [40:0] subW_1119;
wire [66:0] addW_5782;
wire [32:0] slice_1875;
wire [31:0] slice_6538;
wire [50:0] addW_2631;
wire [133:0] concat_7294;
wire [17:0] slice_3387;
wire [33:0] add_4143;
wire [15:0] mul_236;
wire [31:0] slice_4899;
wire [47:0] addW_992;
wire [13:0] slice_5655;
wire [35:0] mul_1748;
wire [19:0] addW_6411;
wire [34:0] addW_2504;
wire [32:0] lsl_7167;
wire [32:0] slice_3260;
wire [27:0] mul_4016;
wire [7:0] slice_109;
wire [7:0] slice_4772;
wire [388:0] addW_865;
wire [8:0] slice_5528;
wire [15:0] slice_1621;
wire [39:0] mul_6284;
wire [50:0] addW_2377;
wire [33:0] add_7040;
wire [35:0] mul_3133;
wire [41:0] subW_3889;
wire [25:0] lsl_4645;
wire [50:0] addW_738;
wire [16:0] mulnw_5401;
wire [17:0] slice_1494;
wire [99:0] addW_6157;
wire [49:0] concat_6913;
wire [7:0] slice_3006;
wire [17:0] slice_3762;
wire [19:0] addW_4518;
wire [15:0] mul_611;
wire [32:0] slice_5274;
wire [65:0] concat_1367;
wire [33:0] addW_6030;
wire [32:0] lsl_2123;
wire [41:0] subW_6786;
wire [26:0] add_2879;
wire [7:0] slice_7542;
wire [133:0] subW_3635;
wire [15:0] mulnw_4391;
wire [32:0] slice_484;
wire [31:0] slice_5147;
wire [65:0] concat_1240;
wire [13:0] slice_5903;
wire [45:0] concat_1996;
wire [16:0] mulnw_6659;
wire [8:0] slice_2752;
wire [7:0] slice_7415;
wire [15:0] slice_3508;
wire [34:0] addW_4264;
wire [49:0] concat_357;
wire [19:0] addW_5020;
wire [35:0] mul_1113;
wire [71:0] subW_5776;
wire [63:0] slice_1869;
wire [39:0] mul_6532;
wire [17:0] add_2625;
wire [17:0] slice_7288;
wire [31:0] slice_3381;
wire [7:0] slice_4137;
wire [7:0] slice_230;
wire [39:0] mul_4893;
wire [45:0] concat_986;
wire [50:0] addW_5649;
wire [13:0] slice_1742;
wire [31:0] mul_6405;
wire [15:0] mulnw_2498;
wire [15:0] mul_7161;
wire [63:0] slice_3254;
wire [17:0] slice_4010;
wire [7:0] slice_103;
wire [8:0] slice_4766;
wire [135:0] subW_859;
wire [33:0] mul_5522;
wire [66:0] concat_1615;
wire [17:0] slice_6278;
wire [17:0] add_2371;
wire [7:0] slice_7034;
wire [13:0] slice_3127;
wire [17:0] slice_3883;
wire [32:0] lsl_4639;
wire [17:0] add_732;
wire [7:0] slice_5395;
wire [31:0] slice_1488;
wire [41:0] subW_6151;
wire [195:0] addW_2244;
wire [16:0] slice_6907;
wire [15:0] slice_3000;
wire [19:0] addW_3756;
wire [27:0] mul_4512;
wire [7:0] slice_605;
wire [34:0] addW_5268;
wire [19:0] addW_1361;
wire [17:0] slice_6024;
wire [31:0] mul_2117;
wire [17:0] slice_6780;
wire [15:0] mulnw_2873;
wire [16:0] mulnw_7536;
wire [70:0] subW_3629;
wire [49:0] concat_4385;
wire [63:0] slice_478;
wire [31:0] slice_5141;
wire [19:0] addW_1234;
wire [127:0] slice_5897;
wire [13:0] slice_1990;
wire [15:0] slice_6653;
wire [17:0] add_2746;
wire [16:0] mulnw_7409;
wire [33:0] addW_3502;
wire [41:0] subW_4258;
wire [16:0] slice_351;
wire [31:0] mul_5014;
wire [15:0] slice_1107;
wire [40:0] subW_5770;
wire [66:0] concat_1863;
wire [17:0] slice_6526;
wire [16:0] mulnw_2619;
wire [19:0] addW_7282;
wire [63:0] slice_3375;
wire [8:0] slice_4131;
wire [15:0] slice_224;
wire [17:0] slice_4887;
wire [13:0] slice_980;
wire [17:0] add_5643;
wire [33:0] add_1736;
wire [31:0] slice_6399;
wire [8:0] slice_2492;
wire [7:0] slice_7155;
wire [66:0] concat_3248;
wire [19:0] addW_4004;
wire [16:0] mulnw_97;
wire [33:0] mul_4760;
wire [70:0] subW_853;
wire [65:0] addW_5516;
wire [15:0] mul_1609;
wire [31:0] slice_6272;
wire [16:0] mulnw_2365;
wire [8:0] slice_7028;
wire [33:0] add_3121;
wire [34:0] addW_3877;
wire [15:0] mul_4633;
wire [16:0] mulnw_726;
wire [15:0] slice_5389;
wire [70:0] subW_1482;
wire [17:0] slice_6145;
wire [71:0] subW_2238;
wire [195:0] concat_6901;
wire [32:0] slice_2994;
wire [27:0] mul_3750;
wire [17:0] slice_4506;
wire [26:0] add_599;
wire [15:0] mulnw_5262;
wire [17:0] slice_1355;
wire [19:0] addW_6018;
wire [16:0] slice_2111;
wire [31:0] slice_6774;
wire [49:0] concat_2867;
wire [7:0] slice_7530;
wire [39:0] mul_3623;
wire [16:0] slice_4379;
wire [66:0] concat_472;
wire [51:0] addW_5135;
wire [17:0] slice_1228;
wire [197:0] addW_5891;
wire [63:0] slice_1984;
wire [32:0] slice_6647;
wire [16:0] mulnw_2740;
wire [7:0] slice_7403;
wire [41:0] subW_3496;
wire [17:0] slice_4252;
wire [65:0] concat_345;
wire [32:0] slice_5008;
wire [47:0] addW_1101;
wire [35:0] mul_5764;
wire [15:0] mul_1857;
wire [13:0] slice_6520;
wire [25:0] lsl_2613;
wire [31:0] mul_7276;
wire [262:0] subW_3369;
wire [33:0] mul_4125;
wire [32:0] slice_218;
wire [31:0] slice_4881;
wire [47:0] addW_974;
wire [16:0] mulnw_5637;
wire [7:0] slice_1730;
wire [39:0] mul_6393;
wire [17:0] add_2486;
wire [15:0] slice_7149;
wire [15:0] mul_3242;
wire [27:0] mul_3998;
wire [16:0] mulnw_91;
wire [32:0] slice_4754;
wire [39:0] mul_847;
wire [68:0] subW_5510;
wire [7:0] slice_1603;
wire [39:0] mul_6266;
wire [25:0] lsl_2359;
wire [33:0] mul_7022;
wire [7:0] slice_3115;
wire [17:0] slice_3871;
wire [7:0] slice_4627;
wire [25:0] lsl_720;
wire [97:0] concat_5383;
wire [39:0] mul_1476;
wire [34:0] addW_6139;
wire [40:0] subW_2232;
wire [67:0] subW_6895;
wire [63:0] slice_2988;
wire [17:0] slice_3744;
wire [19:0] addW_4500;
wire [15:0] mulnw_593;
wire [8:0] slice_5256;
wire [66:0] concat_1349;
wire [27:0] mul_6012;
wire [47:0] addW_2105;
wire [34:0] addW_6768;
wire [16:0] slice_2861;
wire [15:0] slice_7524;
wire [17:0] slice_3617;
wire [195:0] concat_4373;
wire [15:0] mul_466;
wire [49:0] concat_5129;
wire [31:0] slice_1222;
wire [71:0] subW_5885;
wire [134:0] subW_1978;
wire [26:0] add_6641;
wire [15:0] slice_2734;
wire [15:0] slice_7397;
wire [17:0] slice_3490;
wire [31:0] slice_4246;
wire [19:0] addW_339;
wire [26:0] add_5002;
wire [45:0] concat_1095;
wire [15:0] slice_5758;
wire [7:0] slice_1851;
wire [71:0] subW_6514;
wire [32:0] lsl_2607;
wire [32:0] slice_7270;
wire [134:0] subW_3363;
wire [15:0] slice_4119;
wire [26:0] add_4875;
wire [45:0] concat_968;
wire [25:0] lsl_5631;
wire [7:0] slice_1724;
wire [17:0] slice_6387;
wire [16:0] mulnw_2480;
wire [33:0] addW_7143;
wire [7:0] slice_3236;
wire [63:0] slice_3992;
wire [15:0] slice_85;
wire [63:0] slice_4748;
wire [17:0] slice_841;
wire [33:0] add_5504;
wire [26:0] add_1597;
wire [17:0] slice_6260;
wire [32:0] lsl_2353;
wire [32:0] slice_7016;
wire [7:0] slice_3109;
wire [19:0] addW_3865;
wire [15:0] slice_4621;
wire [32:0] lsl_714;
wire [40:0] subW_5377;
wire [17:0] slice_1470;
wire [17:0] slice_6133;
wire [35:0] mul_2226;
wire [26:0] add_6889;
wire [66:0] concat_2982;
wire [19:0] addW_3738;
wire [27:0] mul_4494;
wire [49:0] concat_587;
wire [17:0] add_5250;
wire [15:0] mul_1343;
wire [17:0] slice_6006;
wire [45:0] concat_2099;
wire [15:0] mulnw_6762;
wire [65:0] concat_2855;
wire [66:0] concat_7518;
wire [34:0] addW_3611;
wire [67:0] subW_4367;
wire [7:0] slice_460;
wire [15:0] slice_5123;
wire [67:0] subW_1216;
wire [40:0] subW_5879;
wire [69:0] concat_1972;
wire [16:0] mulnw_6635;
wire [16:0] slice_2728;
wire [32:0] slice_7391;
wire [31:0] slice_3484;
wire [34:0] addW_4240;
wire [17:0] slice_333;
wire [16:0] mulnw_4996;
wire [13:0] slice_1089;
wire [47:0] addW_5752;
wire [26:0] add_1845;
wire [40:0] subW_6508;
wire [31:0] mul_2601;
wire [26:0] add_7264;
wire [69:0] concat_3357;
wire [25:0] lsl_4113;
wire [68:0] subW_206;
wire [16:0] mulnw_4869;
wire [13:0] slice_962;
wire [32:0] lsl_5625;
wire [16:0] mulnw_1718;
wire [31:0] slice_6381;
wire [15:0] slice_2474;
wire [17:0] slice_7137;
wire [26:0] add_3230;
wire [69:0] concat_3986;
wire [16:0] slice_79;
wire [99:0] addW_4742;
wire [34:0] addW_835;
wire [7:0] slice_5498;
wire [15:0] mulnw_1591;
wire [13:0] slice_6254;
wire [31:0] mul_2347;
wire [135:0] subW_7010;
wire [16:0] mulnw_3103;
wire [27:0] mul_3859;
wire [33:0] addW_4615;
wire [31:0] mul_708;
wire [35:0] mul_5371;
wire [34:0] addW_1464;
wire [19:0] addW_6127;
wire [15:0] slice_2220;
wire [16:0] mulnw_6883;
wire [15:0] mul_2976;
wire [27:0] mul_3732;
wire [31:0] slice_4488;
wire [16:0] slice_581;
wire [16:0] mulnw_5244;
wire [7:0] slice_1337;
wire [19:0] addW_6000;
wire [13:0] slice_2093;
wire [8:0] slice_6756;
wire [19:0] addW_2849;
wire [15:0] mul_7512;
wire [41:0] subW_3605;
wire [26:0] add_4361;
wire [26:0] add_454;
wire [65:0] concat_5117;
wire [26:0] add_1210;
wire [35:0] mul_5873;
wire [19:0] addW_1966;
wire [33:0] add_6629;
wire [31:0] slice_2722;
wire [70:0] subW_7385;
wire [41:0] subW_3478;
wire [15:0] mulnw_4234;
wire [65:0] concat_327;
wire [33:0] add_4990;
wire [50:0] addW_1083;
wire [45:0] concat_5746;
wire [15:0] mulnw_1839;
wire [35:0] mul_6502;
wire [16:0] slice_2595;
wire [16:0] mulnw_7258;
wire [19:0] addW_3351;
wire [32:0] lsl_4107;
wire [33:0] add_200;
wire [33:0] add_4863;
wire [130:0] concat_956;
wire [31:0] mul_5619;
wire [7:0] slice_1712;
wire [26:0] add_6375;
wire [32:0] slice_2468;
wire [19:0] addW_7131;
wire [15:0] mulnw_3224;
wire [19:0] addW_3980;
wire [41:0] subW_4736;
wire [50:0] addW_829;
wire [7:0] slice_5492;
wire [49:0] concat_1585;
wire [68:0] subW_6248;
wire [64:0] slice_2341;
wire [70:0] subW_7004;
wire [7:0] slice_3097;
wire [15:0] slice_3853;
wire [17:0] slice_4609;
wire [16:0] slice_702;
wire [13:0] slice_5365;
wire [41:0] subW_1458;
wire [27:0] mul_6121;
wire [47:0] addW_2214;
wire [33:0] add_6877;
wire [7:0] slice_2970;
wire [63:0] slice_3726;
wire [135:0] subW_4482;
wire [64:0] slice_575;
wire [15:0] slice_5238;
wire [26:0] add_1331;
wire [27:0] mul_5994;
wire [47:0] addW_2087;
wire [17:0] add_6750;
wire [17:0] slice_2843;
wire [7:0] slice_7506;
wire [17:0] slice_3599;
wire [16:0] mulnw_4355;
wire [15:0] mulnw_448;
wire [19:0] addW_5111;
wire [16:0] mulnw_1204;
wire [15:0] slice_5867;
wire [17:0] slice_1960;
wire [7:0] slice_6623;
wire [50:0] addW_2716;
wire [39:0] mul_7379;
wire [17:0] slice_3472;
wire [8:0] slice_4228;
wire [19:0] addW_321;
wire [7:0] slice_4984;
wire [17:0] add_1077;
wire [13:0] slice_5740;
wire [49:0] concat_1833;
wire [15:0] slice_6496;
wire [47:0] addW_2589;
wire [33:0] add_7252;
wire [17:0] slice_3345;
wire [15:0] mul_4101;
wire [7:0] slice_194;
wire [7:0] slice_4857;
wire [15:0] slice_950;
wire [64:0] slice_5613;
wire [15:0] slice_1706;
wire [16:0] mulnw_6369;
wire [26:0] add_2462;
wire [27:0] mul_7125;
wire [49:0] concat_3218;
wire [17:0] slice_3974;
wire [47:0] addW_67;
wire [17:0] slice_4730;
wire [17:0] add_823;
wire [16:0] mulnw_5486;
wire [16:0] slice_1579;
wire [33:0] add_6242;
wire [99:0] addW_2335;
wire [39:0] mul_6998;
wire [15:0] slice_3091;
wire [25:0] lsl_3847;
wire [19:0] addW_4603;
wire [47:0] addW_696;
wire [40:0] subW_5359;
wire [17:0] slice_1452;
wire [15:0] slice_6115;
wire [45:0] concat_2208;
wire [7:0] slice_6871;
wire [26:0] add_2964;
wire [66:0] concat_3720;
wire [70:0] subW_4476;
wire [259:0] concat_569;
wire [16:0] slice_5232;
wire [15:0] mulnw_1325;
wire [63:0] slice_5988;
wire [45:0] concat_2081;
wire [16:0] mulnw_6744;
wire [65:0] concat_2837;
wire [26:0] add_7500;
wire [31:0] slice_3593;
wire [33:0] add_4349;
wire [49:0] concat_442;
wire [17:0] slice_5105;
wire [33:0] add_1198;
wire [50:0] addW_5861;
wire [99:0] concat_1954;
wire [8:0] slice_6617;
wire [17:0] add_2710;
wire [17:0] slice_7373;
wire [31:0] slice_3466;
wire [17:0] add_4222;
wire [17:0] slice_315;
wire [8:0] slice_4978;
wire [16:0] mulnw_1071;
wire [50:0] addW_5734;
wire [16:0] slice_1827;
wire [47:0] addW_6490;
wire [45:0] concat_2583;
wire [7:0] slice_7246;
wire [99:0] concat_3339;
wire [7:0] slice_4095;
wire [7:0] slice_188;
wire [8:0] slice_4851;
wire [25:0] lsl_944;
wire [388:0] concat_5607;
wire [257:0] addW_1700;
wire [33:0] add_6363;
wire [16:0] mulnw_2456;
wire [17:0] slice_7119;
wire [16:0] slice_3212;
wire [98:0] concat_3968;
wire [45:0] concat_61;
wire [34:0] addW_4724;
wire [16:0] mulnw_817;
wire [7:0] slice_5480;
wire [195:0] concat_1573;
wire [7:0] slice_6236;
wire [41:0] subW_2329;
wire [17:0] slice_6992;
wire [16:0] slice_3085;
wire [32:0] lsl_3841;
wire [27:0] mul_4597;
wire [45:0] concat_690;
wire [35:0] mul_5353;
wire [31:0] slice_1446;
wire [25:0] lsl_6109;
wire [13:0] slice_2202;
wire [8:0] slice_6865;
wire [15:0] mulnw_2958;
wire [15:0] mul_3714;
wire [39:0] mul_4470;
wire [31:0] slice_563;
wire [31:0] slice_5226;
wire [49:0] concat_1319;
wire [66:0] concat_5982;
wire [13:0] slice_2075;
wire [15:0] slice_6738;
wire [19:0] addW_2831;
wire [15:0] mulnw_7494;
wire [34:0] addW_3587;
wire [7:0] slice_4343;
wire [16:0] slice_436;
wire [66:0] concat_5099;
wire [7:0] slice_1192;
wire [17:0] add_5855;
wire [33:0] add_1948;
wire [33:0] mul_6611;
wire [16:0] mulnw_2704;
wire [34:0] addW_7367;
wire [31:0] slice_3460;
wire [16:0] mulnw_4216;
wire [13:0] slice_309;
wire [33:0] mul_4972;
wire [25:0] lsl_1065;
wire [17:0] add_5728;
wire [65:0] concat_1821;
wire [45:0] concat_6484;
wire [13:0] slice_2577;
wire [8:0] slice_7240;
wire [33:0] add_3333;
wire [15:0] slice_4089;
wire [16:0] mulnw_182;
wire [33:0] mul_4845;
wire [32:0] lsl_938;
wire [132:0] subW_5601;
wire [7:0] slice_6357;
wire [33:0] add_2450;
wire [19:0] addW_7113;
wire [65:0] concat_3206;
wire [40:0] subW_3962;
wire [13:0] slice_55;
wire [17:0] slice_4718;
wire [25:0] lsl_811;
wire [15:0] slice_5474;
wire [67:0] subW_1567;
wire [7:0] slice_6230;
wire [17:0] slice_2323;
wire [34:0] addW_6986;
wire [259:0] concat_3079;
wire [15:0] mul_3835;
wire [17:0] slice_4591;
wire [13:0] slice_684;
wire [63:0] slice_5347;
wire [34:0] addW_1440;
wire [32:0] lsl_6103;
wire [50:0] addW_2196;
wire [33:0] mul_6859;
wire [49:0] concat_2952;
wire [7:0] slice_3708;
wire [17:0] slice_4464;
wire [51:0] addW_557;
wire [50:0] addW_5220;
wire [16:0] slice_1313;
wire [15:0] mul_5976;
wire [130:0] concat_2069;
wire [128:0] slice_6732;
wire [17:0] slice_2825;
wire [49:0] concat_7488;
wire [15:0] mulnw_3581;
wire [8:0] slice_4337;
wire [65:0] concat_430;
wire [15:0] mul_5093;
wire [8:0] slice_1186;
wire [16:0] mulnw_5849;
wire [7:0] slice_1942;
wire [66:0] addW_6605;
wire [25:0] lsl_2698;
wire [41:0] subW_7361;
wire [50:0] addW_3454;
wire [15:0] slice_4210;
wire [195:0] addW_303;
wire [15:0] slice_4966;
wire [32:0] lsl_1059;
wire [16:0] mulnw_5722;
wire [19:0] addW_1815;
wire [13:0] slice_6478;
wire [47:0] addW_2571;
wire [33:0] mul_7234;
wire [7:0] slice_3327;
wire [32:0] slice_4083;
wire [7:0] slice_176;
wire [64:0] slice_4839;
wire [15:0] mul_932;
wire [69:0] concat_5595;
wire [388:0] addW_1688;
wire [8:0] slice_6351;
wire [7:0] slice_2444;
wire [27:0] mul_7107;
wire [19:0] addW_3200;
wire [35:0] mul_3956;
wire [47:0] addW_49;
wire [19:0] addW_4712;
wire [32:0] lsl_805;
wire [97:0] concat_5468;
wire [26:0] add_1561;
wire [16:0] mulnw_6224;
wire [34:0] addW_2317;
wire [34:0] addW_6980;
wire [31:0] slice_3073;
wire [7:0] slice_3829;
wire [19:0] addW_4585;
wire [47:0] addW_678;
wire [260:0] concat_5341;
wire [15:0] mulnw_1434;
wire [15:0] mul_6097;
wire [17:0] add_2190;
wire [31:0] slice_6853;
wire [16:0] slice_2946;
wire [26:0] add_3702;
wire [34:0] addW_4458;
wire [49:0] concat_551;
wire [17:0] add_5214;
wire [194:0] concat_1307;
wire [7:0] slice_5970;
wire [15:0] slice_2063;
wire [258:0] addW_6726;
wire [13:0] slice_2819;
wire [16:0] slice_7482;
wire [8:0] slice_3575;
wire [33:0] mul_4331;
wire [19:0] addW_424;
wire [7:0] slice_5087;
wire [33:0] mul_1180;
wire [25:0] lsl_5843;
wire [7:0] slice_1936;
wire [68:0] subW_6599;
wire [32:0] lsl_2692;
wire [17:0] slice_7355;
wire [17:0] add_3448;
wire [128:0] slice_4204;
wire [71:0] subW_297;
wire [25:0] lsl_4960;
wire [31:0] mul_1053;
wire [25:0] lsl_5716;
wire [17:0] slice_1809;
wire [50:0] addW_6472;
wire [45:0] concat_2565;
wire [15:0] slice_7228;
wire [7:0] slice_3321;
wire [63:0] slice_4077;
wire [15:0] slice_170;
wire [69:0] concat_4833;
wire [7:0] slice_926;
wire [19:0] addW_5589;
wire [135:0] subW_1682;
wire [33:0] mul_6345;
wire [8:0] slice_2438;
wire [63:0] slice_7101;
wire [17:0] slice_3194;
wire [13:0] slice_3950;
wire [27:0] mul_4706;
wire [31:0] mul_799;
wire [40:0] subW_5462;
wire [16:0] mulnw_1555;
wire [7:0] slice_6218;
wire [17:0] slice_2311;
wire [15:0] mulnw_6974;
wire [51:0] addW_3067;
wire [15:0] slice_3823;
wire [27:0] mul_4579;
wire [45:0] concat_672;
wire [32:0] slice_5335;
wire [8:0] slice_1428;
wire [7:0] slice_6091;
wire [16:0] mulnw_2184;
wire [39:0] mul_6847;
wire [65:0] concat_2940;
wire [2054:0] concat_7603;
wire [15:0] mulnw_3696;
wire [34:0] addW_4452;
wire [15:0] slice_545;
wire [16:0] mulnw_5208;
wire [67:0] subW_1301;
wire [26:0] add_5964;
wire [25:0] lsl_2057;
wire [127:0] slice_6720;
wire [195:0] addW_2813;
wire [196:0] concat_7476;
wire [17:0] add_3569;
wire [31:0] slice_4325;
wire [17:0] slice_418;
wire [26:0] add_5081;
wire [31:0] slice_1174;
wire [32:0] lsl_5837;
wire [16:0] mulnw_1930;
wire [33:0] add_6593;
wire [31:0] mul_2686;
wire [31:0] slice_7349;
wire [16:0] mulnw_3442;
wire [257:0] addW_4198;
wire [40:0] subW_291;
wire [32:0] lsl_4954;
wire [65:0] addW_1047;
wire [32:0] lsl_5710;
wire [65:0] concat_1803;
wire [17:0] add_6466;
wire [13:0] slice_2559;
wire [25:0] lsl_7222;
wire [16:0] mulnw_3315;
wire [66:0] concat_4071;
wire [97:0] concat_164;
wire [19:0] addW_4827;
wire [15:0] slice_920;
wire [17:0] slice_5583;
wire [70:0] subW_1676;
wire [65:0] addW_6339;
wire [33:0] mul_2432;
wire [69:0] concat_7095;
wire [65:0] concat_3188;
wire [33:0] add_3944;
wire [17:0] slice_37;
wire [15:0] slice_4700;
wire [16:0] slice_793;
wire [35:0] mul_5456;
wire [33:0] add_1549;
wire [15:0] slice_6212;
wire [19:0] addW_2305;
wire [8:0] slice_6968;
wire [49:0] concat_3061;
wire [32:0] slice_3817;
wire [63:0] slice_4573;
wire [13:0] slice_666;
wire [51:0] addW_5329;
wire [17:0] add_1422;
wire [15:0] slice_6085;
wire [25:0] lsl_2178;
wire [17:0] slice_6841;
wire [19:0] addW_2934;
wire [255:0] slice_7597;
wire [49:0] concat_3690;
wire [15:0] mulnw_4446;
wire [65:0] concat_539;
wire [25:0] lsl_5202;
wire [26:0] add_1295;
wire [15:0] mulnw_5958;
wire [32:0] lsl_2051;
wire [196:0] addW_6714;
wire [71:0] subW_2807;
wire [70:0] subW_7470;
wire [16:0] mulnw_3563;
wire [39:0] mul_4319;
wire [65:0] concat_412;
wire [15:0] mulnw_5075;
wire [39:0] mul_1168;
wire [31:0] mul_5831;
wire [7:0] slice_1924;
wire [7:0] slice_6587;
wire [16:0] slice_2680;
wire [34:0] addW_7343;
wire [25:0] lsl_3436;
wire [262:0] subW_4192;
wire [35:0] mul_285;
wire [15:0] mul_4948;
wire [130:0] concat_1041;
wire [31:0] mul_5704;
wire [19:0] addW_1797;
wire [16:0] mulnw_6460;
wire [13:0] slice_2553;
wire [32:0] lsl_7216;
wire [7:0] slice_3309;
wire [15:0] mul_4065;
wire [40:0] subW_158;
wire [17:0] slice_4821;
wire [33:0] addW_914;
wire [98:0] concat_5577;
wire [39:0] mul_1670;
wire [68:0] subW_6333;
wire [66:0] addW_2426;
wire [19:0] addW_7089;
wire [19:0] addW_3182;
wire [7:0] slice_3938;
wire [31:0] slice_31;
wire [25:0] lsl_4694;
wire [33:0] add_787;
wire [13:0] slice_5450;
wire [7:0] slice_1543;
wire [97:0] concat_6206;
wire [27:0] mul_2299;
wire [17:0] add_6962;
wire [15:0] slice_3055;
wire [63:0] slice_3811;
wire [66:0] concat_4567;
wire [131:0] concat_660;
wire [49:0] concat_5323;
wire [16:0] mulnw_1416;
wire [32:0] slice_6079;
wire [32:0] lsl_2172;
wire [31:0] slice_6835;
wire [17:0] slice_2928;
wire [390:0] addW_7591;
wire [16:0] slice_3684;
wire [8:0] slice_4440;
wire [19:0] addW_533;
wire [32:0] lsl_5196;
wire [16:0] mulnw_1289;
wire [49:0] concat_5952;
wire [15:0] mul_2045;
wire [71:0] subW_6708;
wire [40:0] subW_2801;
wire [39:0] mul_7464;
wire [15:0] slice_3557;
wire [17:0] slice_4313;
wire [19:0] addW_406;
wire [49:0] concat_5069;
wire [17:0] slice_1162;
wire [16:0] slice_5825;
wire [15:0] slice_1918;
wire [7:0] slice_6581;
wire [47:0] addW_2674;
wire [15:0] mulnw_7337;
wire [32:0] lsl_3430;
wire [134:0] subW_4186;
wire [15:0] slice_279;
wire [7:0] slice_4942;
wire [15:0] slice_1035;
wire [64:0] slice_5698;
wire [17:0] slice_1791;
wire [25:0] lsl_6454;
wire [1029:0] concat_2547;
wire [15:0] mul_7210;
wire [15:0] slice_3303;
wire [7:0] slice_4059;
wire [35:0] mul_152;
wire [98:0] concat_4815;
wire [17:0] slice_908;
wire [40:0] subW_5571;
wire [17:0] slice_1664;
wire [33:0] add_6327;
wire [99:0] addW_2420;
wire [17:0] slice_7083;
wire [17:0] slice_3176;
wire [7:0] slice_3932;
wire [13:0] slice_25;
wire [32:0] lsl_4688;
wire [7:0] slice_781;
wire [40:0] subW_5444;
wire [8:0] slice_1537;
wire [40:0] subW_6200;
wire [15:0] slice_2293;
wire [16:0] mulnw_6956;
wire [65:0] concat_3049;
wire [66:0] concat_3805;
wire [15:0] mul_4561;
wire [17:0] slice_654;
wire [15:0] slice_5317;
wire [15:0] slice_1410;
wire [63:0] slice_6073;
wire [31:0] mul_2166;
wire [39:0] mul_6829;
wire [65:0] concat_2922;
wire [135:0] subW_7585;
wire [65:0] concat_3678;
wire [17:0] add_4434;
wire [17:0] slice_527;
wire [31:0] mul_5190;
wire [33:0] add_1283;
wire [16:0] slice_5946;
wire [7:0] slice_2039;
wire [40:0] subW_6702;
wire [35:0] mul_2795;
wire [17:0] slice_7458;
wire [16:0] slice_3551;
wire [31:0] slice_4307;
wire [17:0] slice_400;
wire [16:0] slice_5063;
wire [31:0] slice_1156;
wire [33:0] add_5819;
wire [66:0] concat_1912;
wire [16:0] mulnw_6575;
wire [45:0] concat_2668;
wire [8:0] slice_7331;
wire [31:0] mul_3424;
wire [69:0] concat_4180;
wire [65:0] concat_273;
wire [15:0] slice_4936;
wire [25:0] lsl_1029;
wire [99:0] addW_5692;
wire [31:0] slice_1785;
wire [32:0] lsl_6448;
wire [127:0] slice_2541;
wire [7:0] slice_7204;
wire [66:0] concat_3297;
wire [26:0] add_4053;
wire [13:0] slice_146;
wire [40:0] subW_4809;
wire [19:0] addW_902;
wire [35:0] mul_5565;
wire [34:0] addW_1658;
wire [7:0] slice_6321;
wire [41:0] subW_2414;
wire [98:0] concat_7077;
wire [31:0] slice_3170;
wire [16:0] mulnw_3926;
wire [63:0] slice_19;
wire [15:0] mul_4682;
wire [7:0] slice_775;
wire [35:0] mul_5438;
wire [33:0] mul_1531;
wire [35:0] mul_6194;
wire [25:0] lsl_2287;
wire [15:0] slice_6950;
wire [19:0] addW_3043;
wire [15:0] mul_3799;
wire [7:0] slice_4555;
wire [19:0] addW_648;
wire [66:0] concat_5311;
wire [129:0] addW_1404;
wire [66:0] concat_6067;
wire [65:0] addW_2160;
wire [17:0] slice_6823;
wire [19:0] addW_2916;
wire [70:0] subW_7579;
wire [19:0] addW_3672;
wire [16:0] mulnw_4428;
wire [66:0] concat_521;
wire [16:0] slice_5184;
wire [7:0] slice_1277;
wire [65:0] concat_5940;
wire [15:0] slice_2033;
wire [35:0] mul_6696;
wire [15:0] slice_2789;
wire [34:0] addW_7452;
wire [31:0] slice_3545;
wire [39:0] mul_4301;
wire [31:0] slice_394;
wire [16:0] slice_5057;
wire [39:0] mul_1150;
wire [7:0] slice_5813;
wire [15:0] mul_1906;
wire [7:0] slice_6569;
wire [13:0] slice_2662;
wire [17:0] add_7325;
wire [16:0] slice_3418;
wire [19:0] addW_4174;
wire [19:0] addW_267;
wire [32:0] slice_4930;
wire [32:0] lsl_1023;
wire [41:0] subW_5686;
wire [70:0] subW_1779;
wire [31:0] mul_6442;
wire [197:0] addW_2535;
wire [15:0] slice_7198;
wire [15:0] mul_3291;
wire [15:0] mulnw_4047;
wire [40:0] subW_140;
wire [35:0] mul_4803;
wire [27:0] mul_896;
wire [13:0] slice_5559;
wire [34:0] addW_1652;
wire [7:0] slice_6315;
wire [17:0] slice_2408;
wire [40:0] subW_7071;
wire [70:0] subW_3164;
wire [7:0] slice_3920;
wire [255:0] slice_13;
wire [7:0] slice_4676;
wire [16:0] mulnw_769;
wire [63:0] slice_5432;
wire [31:0] slice_1525;
wire [13:0] slice_6188;
wire [32:0] lsl_2281;
wire [32:0] slice_6944;
wire [17:0] slice_3037;
wire [7:0] slice_3793;
wire [26:0] add_4549;
wire [31:0] mul_642;
wire [15:0] mul_5305;
wire [127:0] slice_1398;
wire [15:0] mul_6061;
wire [130:0] concat_2154;
wire [13:0] slice_6817;
wire [17:0] slice_2910;
wire [39:0] mul_7573;
wire [17:0] slice_3666;
wire [15:0] slice_4422;
wire [15:0] mul_515;
wire [47:0] addW_5178;
wire [8:0] slice_1271;
wire [19:0] addW_5934;
wire [33:0] addW_2027;
wire [15:0] slice_6690;
wire [47:0] addW_2783;
wire [41:0] subW_7446;
wire [50:0] addW_3539;
wire [17:0] slice_4295;
wire [67:0] subW_388;
wire [17:0] slice_1144;
wire [7:0] slice_5807;
wire [7:0] slice_1900;
wire [15:0] slice_6563;
wire [47:0] addW_2656;
wire [16:0] mulnw_7319;
wire [47:0] addW_3412;
wire [17:0] slice_4168;
wire [17:0] slice_261;
wire [64:0] slice_4924;
wire [15:0] mul_1017;
wire [17:0] slice_5680;
wire [39:0] mul_1773;
wire [64:0] slice_6436;
wire [71:0] subW_2529;
wire [32:0] slice_7192;
wire [7:0] slice_3285;
wire [49:0] concat_4041;
wire [35:0] mul_134;
wire [13:0] slice_4797;
wire [17:0] slice_890;
wire [33:0] add_5553;
wire [15:0] mulnw_1646;
wire [16:0] mulnw_6309;
wire [34:0] addW_2402;
wire [35:0] mul_7065;
wire [39:0] mul_3158;
wire [15:0] slice_3914;
wire [15:0] slice_4670;
wire [7:0] slice_763;
wire [98:0] addW_5426;
wire [39:0] mul_1519;
wire [40:0] subW_6182;
wire [15:0] mul_2275;
wire [26:0] add_6938;
wire [66:0] concat_3031;
wire [26:0] add_3787;
wire [15:0] mulnw_4543;
wire [31:0] slice_636;
wire [7:0] slice_5299;
wire [131:0] concat_1392;
wire [7:0] slice_6055;
wire [15:0] slice_2148;
wire [71:0] subW_6811;
wire [31:0] slice_2904;
wire [17:0] slice_7567;
wire [65:0] concat_3660;
wire [32:0] slice_4416;
wire [7:0] slice_509;
wire [45:0] concat_5172;
wire [33:0] mul_1265;
wire [17:0] slice_5928;
wire [17:0] slice_2021;
wire [50:0] addW_6684;
wire [45:0] concat_2777;
wire [17:0] slice_7440;
wire [17:0] add_3533;
wire [13:0] slice_4289;
wire [26:0] add_382;
wire [773:0] addW_5045;
wire [127:0] slice_1138;
wire [16:0] mulnw_5801;
wire [26:0] add_1894;
wire [97:0] concat_6557;
wire [45:0] concat_2650;
wire [15:0] slice_7313;
wire [45:0] concat_3406;
wire [99:0] concat_4162;
wire [66:0] concat_255;
wire [69:0] concat_4918;
wire [7:0] slice_1011;
wire [34:0] addW_5674;
wire [17:0] slice_1767;
wire [387:0] concat_6430;
wire [40:0] subW_2523;
wire [63:0] slice_7186;
wire [26:0] add_3279;
wire [16:0] slice_4035;
wire [63:0] slice_128;
wire [33:0] add_4791;
wire [19:0] addW_884;
wire [7:0] slice_5547;
wire [8:0] slice_1640;
wire [7:0] slice_6303;
wire [17:0] slice_2396;
wire [13:0] slice_7059;
wire [17:0] slice_3152;
wire [16:0] slice_3908;
wire [32:0] slice_4664;
wire [15:0] slice_757;
wire [34:0] addW_5420;
wire [17:0] slice_1513;
wire [35:0] mul_6176;
wire [7:0] slice_2269;
wire [16:0] mulnw_6932;
wire [15:0] mul_3025;
wire [15:0] mulnw_3781;
wire [49:0] concat_4537;
wire [39:0] mul_630;
wire [26:0] add_5293;
wire [17:0] slice_1386;
wire [26:0] add_6049;
wire [25:0] lsl_2142;
wire [40:0] subW_6805;
wire [67:0] subW_2898;
wire [34:0] addW_7561;
wire [19:0] addW_3654;
wire [26:0] add_4410;
wire [26:0] add_503;
wire [13:0] slice_5166;
wire [31:0] slice_1259;
wire [65:0] concat_5922;
wire [19:0] addW_2015;
wire [17:0] add_6678;
wire [13:0] slice_2771;
wire [31:0] slice_7434;
wire [16:0] mulnw_3527;
wire [71:0] subW_4283;
wire [16:0] mulnw_376;
wire [264:0] subW_5039;
wire [63:0] slice_1132;
wire [7:0] slice_5795;
wire [15:0] mulnw_1888;
wire [40:0] subW_6551;
wire [13:0] slice_2644;
wire [130:0] addW_7307;
wire [13:0] slice_3400;
wire [33:0] add_4156;
wire [15:0] mul_249;
wire [19:0] addW_4912;
wire [15:0] slice_1005;
wire [17:0] slice_5668;
wire [34:0] addW_1761;
wire [132:0] subW_6424;
wire [35:0] mul_2517;
wire [66:0] concat_7180;
wire [15:0] mulnw_3273;
wire [65:0] concat_4029;
wire [98:0] addW_122;
wire [7:0] slice_4785;
wire [27:0] mul_878;
wire [7:0] slice_5541;
wire [17:0] add_1634;
wire [15:0] slice_6297;
wire [19:0] addW_2390;
wire [33:0] add_7053;
wire [34:0] addW_3146;
wire [259:0] concat_3902;
wire [63:0] slice_4658;
wire [32:0] slice_751;
wire [15:0] mulnw_5414;
wire [31:0] slice_1507;
wire [63:0] slice_6170;
wire [15:0] slice_2263;
wire [33:0] add_6926;
wire [7:0] slice_3019;
wire [49:0] concat_3775;
wire [16:0] slice_4531;
wire [17:0] slice_624;
wire [15:0] mulnw_5287;
wire [19:0] addW_1380;
wire [15:0] mulnw_6043;
wire [32:0] lsl_2136;
wire [35:0] mul_6799;
wire [26:0] add_2892;
wire [34:0] addW_7555;
wire [17:0] slice_3648;
wire [16:0] mulnw_4404;
wire [15:0] mulnw_497;
wire [47:0] addW_5160;
wire [39:0] mul_1253;
wire [19:0] addW_5916;
wire [27:0] mul_2009;
wire [16:0] mulnw_6672;
wire [50:0] addW_2765;
wire [34:0] addW_7428;
wire [25:0] lsl_3521;
wire [40:0] subW_4277;
wire [33:0] add_370;
wire [134:0] subW_5033;
wire [99:0] addW_1126;
wire [15:0] slice_5789;
wire [49:0] concat_1882;
wire [35:0] mul_6545;
wire [130:0] concat_2638;
wire [389:0] concat_7301;
wire [47:0] addW_3394;
wire [7:0] slice_4150;
wire [7:0] slice_243;
wire [17:0] slice_4906;
wire [33:0] addW_999;
wire [19:0] addW_5662;
wire [41:0] subW_1755;
wire [69:0] concat_6418;
wire [15:0] slice_2511;
wire [15:0] mul_7174;
wire [49:0] concat_3267;
wire [19:0] addW_4023;
wire [34:0] addW_116;
wire [7:0] slice_4779;
wire [13:0] slice_872;
wire [16:0] mulnw_5535;
wire [16:0] mulnw_1628;
wire [97:0] concat_6291;
wire [27:0] mul_2384;
wire [7:0] slice_7047;
wire [41:0] subW_3140;
wire [31:0] slice_3896;
wire [66:0] concat_4652;
wire [130:0] concat_745;
wire [8:0] slice_5408;
wire [39:0] mul_1501;
wire [259:0] concat_6164;
wire [32:0] slice_2257;
wire [7:0] slice_6920;
wire [26:0] add_3013;
wire [16:0] slice_3769;
wire [65:0] concat_4525;
wire [31:0] slice_618;
wire [49:0] concat_5281;
wire [31:0] mul_1374;
wire [49:0] concat_6037;
wire [15:0] mul_2130;
wire [15:0] slice_6793;
wire [16:0] mulnw_2886;
wire [15:0] mulnw_7549;
wire [13:0] slice_3642;
wire [33:0] add_4398;
wire [49:0] concat_491;
wire [45:0] concat_5154;
wire [17:0] slice_1247;
wire [17:0] slice_5910;
wire [17:0] slice_2003;
wire [25:0] lsl_6666;
wire [17:0] add_2759;
wire [15:0] mulnw_7422;
wire [32:0] lsl_3515;
wire [35:0] mul_4271;
wire [7:0] slice_364;
wire [69:0] concat_5027;
wire [41:0] subW_1120;
wire [32:0] slice_5783;
wire [16:0] slice_1876;
wire [13:0] slice_6539;
wire [15:0] slice_2632;
wire [134:0] subW_7295;
wire [45:0] concat_3388;
wire [7:0] slice_4144;
wire [26:0] add_237;
wire [98:0] concat_4900;
wire [17:0] slice_993;
wire [27:0] mul_5656;
wire [17:0] slice_1749;
wire [19:0] addW_6412;
wire [50:0] addW_2505;
wire [7:0] slice_7168;
wire [16:0] slice_3261;
wire [17:0] slice_4017;
wire [15:0] mulnw_110;
wire [16:0] mulnw_4773;
wire [127:0] slice_866;
wire [7:0] slice_5529;
wire [15:0] slice_1622;
wire [40:0] subW_6285;
wire [15:0] slice_2378;
wire [7:0] slice_7041;
wire [17:0] slice_3134;
wire [51:0] addW_3890;
wire [15:0] mul_4646;
wire [15:0] slice_739;
wire [17:0] add_5402;
wire [17:0] slice_1495;
wire [31:0] slice_6158;
wire [130:0] addW_2251;
wire [8:0] slice_6914;
wire [15:0] mulnw_3007;
wire [65:0] concat_3763;
wire [19:0] addW_4519;
wire [26:0] add_612;
wire [16:0] slice_5275;
wire [31:0] slice_1368;
wire [16:0] slice_6031;
wire [7:0] slice_2124;
wire [47:0] addW_6787;
wire [33:0] add_2880;
wire [8:0] slice_7543;
wire [195:0] addW_3636;
wire [7:0] slice_4392;
wire [16:0] slice_485;
wire [13:0] slice_5148;
wire [31:0] slice_1241;
wire [255:0] slice_5904;
wire [19:0] addW_1997;
wire [32:0] lsl_6660;
wire [16:0] mulnw_2753;
wire [8:0] slice_7416;
wire [31:0] mul_3509;
wire [15:0] slice_4265;
wire [8:0] slice_358;
wire [19:0] addW_5021;
wire [17:0] slice_1114;
wire [99:0] addW_5777;
wire [195:0] concat_1870;
wire [40:0] subW_6533;
wire [25:0] lsl_2626;
wire [69:0] concat_7289;
wire [13:0] slice_3382;
wire [16:0] mulnw_4138;
wire [15:0] mulnw_231;
wire [40:0] subW_4894;
wire [19:0] addW_987;
wire [15:0] slice_5650;
wire [31:0] slice_1743;
wire [17:0] slice_6406;
wire [17:0] add_2499;
wire [26:0] add_7162;
wire [195:0] concat_3255;
wire [65:0] concat_4011;
wire [8:0] slice_104;
wire [7:0] slice_4767;
wire [196:0] addW_860;
wire [15:0] slice_5523;
wire [32:0] slice_1616;
wire [35:0] mul_6279;
wire [25:0] lsl_2372;
wire [16:0] mulnw_7035;
wire [31:0] slice_3128;
wire [49:0] concat_3884;
wire [7:0] slice_4640;
wire [25:0] lsl_733;
wire [16:0] mulnw_5396;
wire [13:0] slice_1489;
wire [51:0] addW_6152;
wire [63:0] slice_2245;
wire [33:0] mul_6908;
wire [49:0] concat_3001;
wire [19:0] addW_3757;
wire [17:0] slice_4513;
wire [16:0] mulnw_606;
wire [50:0] addW_5269;
wire [39:0] mul_1362;
wire [65:0] concat_6025;
wire [15:0] slice_2118;
wire [45:0] concat_6781;
wire [7:0] slice_2874;
wire [17:0] add_7537;
wire [71:0] subW_3630;
wire [8:0] slice_4386;
wire [194:0] concat_479;
wire [131:0] concat_5142;
wire [39:0] mul_1235;
wire [517:0] concat_5898;
wire [27:0] mul_1991;
wire [31:0] mul_6654;
wire [25:0] lsl_2747;
wire [17:0] add_7410;
wire [16:0] slice_3503;
wire [47:0] addW_4259;
wire [33:0] mul_352;
wire [17:0] slice_5015;
wire [34:0] addW_1108;
wire [41:0] subW_5771;
wire [67:0] subW_1864;
wire [35:0] mul_6527;
wire [32:0] lsl_2620;
wire [19:0] addW_7283;
wire [31:0] slice_3376;
wire [7:0] slice_4132;
wire [49:0] concat_225;
wire [35:0] mul_4888;
wire [27:0] mul_981;
wire [25:0] lsl_5644;
wire [34:0] addW_1737;
wire [98:0] concat_6400;
wire [16:0] mulnw_2493;
wire [15:0] mulnw_7156;
wire [67:0] subW_3249;
wire [19:0] addW_4005;
wire [17:0] add_98;
wire [15:0] slice_4761;
wire [71:0] subW_854;
wire [32:0] slice_5517;
wire [26:0] add_1610;
wire [13:0] slice_6273;
wire [32:0] lsl_2366;
wire [7:0] slice_7029;
wire [34:0] addW_3122;
wire [15:0] slice_3878;
wire [26:0] add_4634;
wire [32:0] lsl_727;
wire [15:0] slice_5390;
wire [71:0] subW_1483;
wire [49:0] concat_6146;
wire [99:0] addW_2239;
wire [66:0] addW_6902;
wire [16:0] slice_2995;
wire [17:0] slice_3751;
wire [65:0] concat_4507;
wire [33:0] add_600;
wire [17:0] add_5263;
wire [17:0] slice_1356;
wire [19:0] addW_6019;
wire [33:0] addW_2112;
wire [13:0] slice_6775;
wire [8:0] slice_2868;
wire [16:0] mulnw_7531;
wire [40:0] subW_3624;
wire [33:0] mul_4380;
wire [67:0] subW_473;
wire [17:0] slice_5136;
wire [17:0] slice_1229;
wire [64:0] slice_5892;
wire [31:0] slice_1985;
wire [16:0] slice_6648;
wire [32:0] lsl_2741;
wire [16:0] mulnw_7404;
wire [47:0] addW_3497;
wire [45:0] concat_4253;
wire [31:0] slice_346;
wire [99:0] concat_5009;
wire [17:0] slice_1102;
wire [17:0] slice_5765;
wire [26:0] add_1858;
wire [63:0] slice_6521;
wire [15:0] mul_2614;
wire [17:0] slice_7277;
wire [388:0] addW_3370;
wire [15:0] slice_4126;
wire [16:0] slice_219;
wire [13:0] slice_4882;
wire [17:0] slice_975;
wire [32:0] lsl_5638;
wire [15:0] mulnw_1731;
wire [40:0] subW_6394;
wire [25:0] lsl_2487;
wire [49:0] concat_7150;
wire [26:0] add_3243;
wire [17:0] slice_3999;
wire [32:0] lsl_92;
wire [16:0] slice_4755;
wire [40:0] subW_848;
wire [98:0] addW_5511;
wire [16:0] mulnw_1604;
wire [40:0] subW_6267;
wire [15:0] mul_2360;
wire [15:0] slice_7023;
wire [15:0] mulnw_3116;
wire [65:0] concat_3872;
wire [15:0] mulnw_4628;
wire [15:0] mul_721;
wire [33:0] addW_5384;
wire [40:0] subW_1477;
wire [15:0] slice_6140;
wire [41:0] subW_2233;
wire [68:0] subW_6896;
wire [194:0] concat_2989;
wire [65:0] concat_3745;
wire [19:0] addW_4501;
wire [7:0] slice_594;
wire [16:0] mulnw_5257;
wire [31:0] slice_1350;
wire [17:0] slice_6013;
wire [17:0] slice_2106;
wire [50:0] addW_6769;
wire [33:0] mul_2862;
wire [15:0] slice_7525;
wire [35:0] mul_3618;
wire [66:0] addW_4374;
wire [26:0] add_467;
wire [19:0] addW_5130;
wire [13:0] slice_1223;
wire [100:0] addW_5886;
wire [135:0] subW_1979;
wire [33:0] add_6642;
wire [31:0] mul_2735;
wire [15:0] slice_7398;
wire [45:0] concat_3491;
wire [13:0] slice_4247;
wire [39:0] mul_340;
wire [33:0] add_5003;
wire [19:0] addW_1096;
wire [34:0] addW_5759;
wire [16:0] mulnw_1852;
wire [99:0] addW_6515;
wire [7:0] slice_2608;
wire [99:0] concat_7271;
wire [135:0] subW_3364;
wire [66:0] concat_4120;
wire [33:0] add_4876;
wire [19:0] addW_969;
wire [15:0] mul_5632;
wire [8:0] slice_1725;
wire [35:0] mul_6388;
wire [32:0] lsl_2481;
wire [16:0] slice_7144;
wire [16:0] mulnw_3237;
wire [31:0] slice_3993;
wire [49:0] concat_86;
wire [259:0] concat_4749;
wire [35:0] mul_842;
wire [34:0] addW_5505;
wire [33:0] add_1598;
wire [35:0] mul_6261;
wire [7:0] slice_2354;
wire [16:0] slice_7017;
wire [8:0] slice_3110;
wire [19:0] addW_3866;
wire [49:0] concat_4622;
wire [7:0] slice_715;
wire [41:0] subW_5378;
wire [35:0] mul_1471;
wire [65:0] concat_6134;
wire [17:0] slice_2227;
wire [33:0] add_6890;
wire [67:0] subW_2983;
wire [19:0] addW_3739;
wire [17:0] slice_4495;
wire [8:0] slice_588;
wire [25:0] lsl_5251;
wire [26:0] add_1344;
wire [65:0] concat_6007;
wire [19:0] addW_2100;
wire [17:0] add_6763;
wire [31:0] slice_2856;
wire [32:0] slice_7519;
wire [15:0] slice_3612;
wire [68:0] subW_4368;
wire [16:0] mulnw_461;
wire [31:0] mul_5124;
wire [68:0] subW_1217;
wire [41:0] subW_5880;
wire [70:0] subW_1973;
wire [7:0] slice_6636;
wire [65:0] addW_2729;
wire [16:0] slice_7392;
wire [13:0] slice_3485;
wire [50:0] addW_4241;
wire [17:0] slice_334;
wire [7:0] slice_4997;
wire [27:0] mul_1090;
wire [17:0] slice_5753;
wire [33:0] add_1846;
wire [41:0] subW_6509;
wire [15:0] slice_2602;
wire [33:0] add_7265;
wire [70:0] subW_3358;
wire [15:0] mul_4114;
wire [98:0] addW_207;
wire [7:0] slice_4870;
wire [27:0] mul_963;
wire [7:0] slice_5626;
wire [17:0] add_1719;
wire [13:0] slice_6382;
wire [31:0] mul_2475;
wire [65:0] concat_7138;
wire [33:0] add_3231;
wire [70:0] subW_3987;
wire [33:0] mul_80;
wire [31:0] slice_4743;
wire [15:0] slice_836;
wire [15:0] mulnw_5499;
wire [7:0] slice_1592;
wire [63:0] slice_6255;
wire [15:0] slice_2348;
wire [196:0] addW_7011;
wire [17:0] add_3104;
wire [17:0] slice_3860;
wire [16:0] slice_4616;
wire [15:0] slice_709;
wire [17:0] slice_5372;
wire [15:0] slice_1465;
wire [19:0] addW_6128;
wire [34:0] addW_2221;
wire [7:0] slice_6884;
wire [26:0] add_2977;
wire [17:0] slice_3733;
wire [13:0] slice_4489;
wire [33:0] mul_582;
wire [32:0] lsl_5245;
wire [16:0] mulnw_1338;
wire [19:0] addW_6001;
wire [27:0] mul_2094;
wire [16:0] mulnw_6757;
wire [39:0] mul_2850;
wire [26:0] add_7513;
wire [47:0] addW_3606;
wire [33:0] add_4362;
wire [33:0] add_455;
wire [31:0] slice_5118;
wire [33:0] add_1211;
wire [17:0] slice_5874;
wire [39:0] mul_1967;
wire [7:0] slice_6630;
wire [130:0] concat_2723;
wire [71:0] subW_7386;
wire [47:0] addW_3479;
wire [17:0] add_4235;
wire [31:0] slice_328;
wire [7:0] slice_4991;
wire [15:0] slice_1084;
wire [19:0] addW_5747;
wire [7:0] slice_1840;
wire [17:0] slice_6503;
wire [33:0] addW_2596;
wire [7:0] slice_7259;
wire [39:0] mul_3352;
wire [7:0] slice_4108;
wire [34:0] addW_201;
wire [7:0] slice_4864;
wire [63:0] slice_957;
wire [15:0] slice_5620;
wire [16:0] mulnw_1713;
wire [33:0] add_6376;
wire [16:0] slice_2469;
wire [19:0] addW_7132;
wire [7:0] slice_3225;
wire [39:0] mul_3981;
wire [51:0] addW_4737;
wire [15:0] slice_830;
wire [8:0] slice_5493;
wire [8:0] slice_1586;
wire [98:0] addW_6249;
wire [32:0] slice_2342;
wire [71:0] subW_7005;
wire [16:0] mulnw_3098;
wire [66:0] concat_3854;
wire [65:0] concat_4610;
wire [33:0] addW_703;
wire [31:0] slice_5366;
wire [47:0] addW_1459;
wire [17:0] slice_6122;
wire [17:0] slice_2215;
wire [7:0] slice_6878;
wire [16:0] mulnw_2971;
wire [31:0] slice_3727;
wire [196:0] addW_4483;
wire [32:0] slice_576;
wire [31:0] mul_5239;
wire [33:0] add_1332;
wire [17:0] slice_5995;
wire [17:0] slice_2088;
wire [25:0] lsl_6751;
wire [17:0] slice_2844;
wire [16:0] mulnw_7507;
wire [45:0] concat_3600;
wire [7:0] slice_4356;
wire [7:0] slice_449;
wire [39:0] mul_5112;
wire [7:0] slice_1205;
wire [34:0] addW_5868;
wire [17:0] slice_1961;
wire [16:0] mulnw_6624;
wire [15:0] slice_2717;
wire [40:0] subW_7380;
wire [45:0] concat_3473;
wire [16:0] mulnw_4229;
wire [39:0] mul_322;
wire [16:0] mulnw_4985;
wire [25:0] lsl_1078;
wire [27:0] mul_5741;
wire [8:0] slice_1834;
wire [34:0] addW_6497;
wire [17:0] slice_2590;
wire [7:0] slice_7253;
wire [17:0] slice_3346;
wire [26:0] add_4102;
wire [15:0] mulnw_195;
wire [16:0] mulnw_4858;
wire [66:0] concat_951;
wire [32:0] slice_5614;
wire [15:0] slice_1707;
wire [7:0] slice_6370;
wire [33:0] add_2463;
wire [17:0] slice_7126;
wire [8:0] slice_3219;
wire [17:0] slice_3975;
wire [17:0] slice_68;
wire [49:0] concat_4731;
wire [25:0] lsl_824;
wire [17:0] add_5487;
wire [33:0] mul_1580;
wire [34:0] addW_6243;
wire [31:0] slice_2336;
wire [40:0] subW_6999;
wire [15:0] slice_3092;
wire [15:0] mul_3848;
wire [19:0] addW_4604;
wire [17:0] slice_697;
wire [41:0] subW_5360;
wire [45:0] concat_1453;
wire [66:0] concat_6116;
wire [19:0] addW_2209;
wire [16:0] mulnw_6872;
wire [33:0] add_2965;
wire [67:0] subW_3721;
wire [71:0] subW_4477;
wire [127:0] slice_570;
wire [66:0] addW_5233;
wire [7:0] slice_1326;
wire [31:0] slice_5989;
wire [19:0] addW_2082;
wire [32:0] lsl_6745;
wire [31:0] slice_2838;
wire [33:0] add_7501;
wire [13:0] slice_3594;
wire [7:0] slice_4350;
wire [8:0] slice_443;
wire [17:0] slice_5106;
wire [7:0] slice_1199;
wire [15:0] slice_5862;
wire [34:0] addW_1955;
wire [7:0] slice_6618;
wire [25:0] lsl_2711;
wire [35:0] mul_7374;
wire [13:0] slice_3467;
wire [25:0] lsl_4223;
wire [17:0] slice_316;
wire [7:0] slice_4979;
wire [32:0] lsl_1072;
wire [15:0] slice_5735;
wire [33:0] mul_1828;
wire [17:0] slice_6491;
wire [19:0] addW_2584;
wire [16:0] mulnw_7247;
wire [34:0] addW_3340;
wire [15:0] mulnw_4096;
wire [8:0] slice_189;
wire [7:0] slice_4852;
wire [15:0] mul_945;
wire [130:0] addW_5608;
wire [128:0] slice_1701;
wire [7:0] slice_6364;
wire [7:0] slice_2457;
wire [65:0] concat_7120;
wire [33:0] mul_3213;
wire [34:0] addW_3969;
wire [19:0] addW_62;
wire [15:0] slice_4725;
wire [32:0] lsl_818;
wire [16:0] mulnw_5481;
wire [66:0] addW_1574;
wire [15:0] mulnw_6237;
wire [51:0] addW_2330;
wire [35:0] mul_6993;
wire [129:0] addW_3086;
wire [7:0] slice_3842;
wire [17:0] slice_4598;
wire [19:0] addW_691;
wire [17:0] slice_5354;
wire [13:0] slice_1447;
wire [15:0] mul_6110;
wire [27:0] mul_2203;
wire [7:0] slice_6866;
wire [7:0] slice_2959;
wire [26:0] add_3715;
wire [40:0] subW_4471;
wire [131:0] concat_564;
wire [130:0] concat_5227;
wire [8:0] slice_1320;
wire [67:0] subW_5983;
wire [27:0] mul_2076;
wire [31:0] mul_6739;
wire [39:0] mul_2832;
wire [7:0] slice_7495;
wire [50:0] addW_3588;
wire [16:0] mulnw_4344;
wire [33:0] mul_437;
wire [31:0] slice_5100;
wire [16:0] mulnw_1193;
wire [25:0] lsl_5856;
wire [34:0] addW_1949;
wire [15:0] slice_6612;
wire [32:0] lsl_2705;
wire [15:0] slice_7368;
wire [130:0] concat_3461;
wire [32:0] lsl_4217;
wire [127:0] slice_310;
wire [15:0] slice_4973;
wire [15:0] mul_1066;
wire [25:0] lsl_5729;
wire [31:0] slice_1822;
wire [19:0] addW_6485;
wire [27:0] mul_2578;
wire [7:0] slice_7241;
wire [34:0] addW_3334;
wire [49:0] concat_4090;
wire [17:0] add_183;
wire [15:0] slice_4846;
wire [7:0] slice_939;
wire [133:0] subW_5602;
wire [257:0] addW_1695;
wire [16:0] mulnw_6358;
wire [7:0] slice_2451;
wire [19:0] addW_7114;
wire [31:0] slice_3207;
wire [41:0] subW_3963;
wire [27:0] mul_56;
wire [65:0] concat_4719;
wire [15:0] mul_812;
wire [15:0] slice_5475;
wire [68:0] subW_1568;
wire [8:0] slice_6231;
wire [49:0] concat_2324;
wire [15:0] slice_6987;
wire [127:0] slice_3080;
wire [26:0] add_3836;
wire [65:0] concat_4592;
wire [27:0] mul_685;
wire [31:0] slice_5348;
wire [50:0] addW_1441;
wire [7:0] slice_6104;
wire [15:0] slice_2197;
wire [15:0] slice_6860;
wire [8:0] slice_2953;
wire [16:0] mulnw_3709;
wire [35:0] mul_4465;
wire [17:0] slice_558;
wire [15:0] slice_5221;
wire [33:0] mul_1314;
wire [26:0] add_5977;
wire [63:0] slice_2070;
wire [64:0] slice_6733;
wire [17:0] slice_2826;
wire [8:0] slice_7489;
wire [17:0] add_3582;
wire [7:0] slice_4338;
wire [31:0] slice_431;
wire [26:0] add_5094;
wire [7:0] slice_1187;
wire [32:0] lsl_5850;
wire [15:0] mulnw_1943;
wire [32:0] slice_6606;
wire [15:0] mul_2699;
wire [47:0] addW_7362;
wire [15:0] slice_3455;
wire [31:0] mul_4211;
wire [63:0] slice_304;
wire [66:0] concat_4967;
wire [7:0] slice_1060;
wire [32:0] lsl_5723;
wire [39:0] mul_1816;
wire [27:0] mul_6479;
wire [17:0] slice_2572;
wire [15:0] slice_7235;
wire [15:0] mulnw_3328;
wire [16:0] slice_4084;
wire [16:0] mulnw_177;
wire [32:0] slice_4840;
wire [26:0] add_933;
wire [70:0] subW_5596;
wire [127:0] slice_1689;
wire [7:0] slice_6352;
wire [16:0] mulnw_2445;
wire [17:0] slice_7108;
wire [39:0] mul_3201;
wire [17:0] slice_3957;
wire [17:0] slice_50;
wire [19:0] addW_4713;
wire [7:0] slice_806;
wire [33:0] addW_5469;
wire [33:0] add_1562;
wire [17:0] add_6225;
wire [15:0] slice_2318;
wire [50:0] addW_6981;
wire [131:0] concat_3074;
wire [15:0] mulnw_3830;
wire [19:0] addW_4586;
wire [17:0] slice_679;
wire [127:0] slice_5342;
wire [17:0] add_1435;
wire [26:0] add_6098;
wire [25:0] lsl_2191;
wire [97:0] concat_6854;
wire [33:0] mul_2947;
wire [33:0] add_3703;
wire [15:0] slice_4459;
wire [19:0] addW_552;
wire [25:0] lsl_5215;
wire [65:0] addW_1308;
wire [16:0] mulnw_5971;
wire [66:0] concat_2064;
wire [128:0] slice_6727;
wire [127:0] slice_2820;
wire [33:0] mul_7483;
wire [16:0] mulnw_3576;
wire [15:0] slice_4332;
wire [39:0] mul_425;
wire [16:0] mulnw_5088;
wire [15:0] slice_1181;
wire [15:0] mul_5844;
wire [8:0] slice_1937;
wire [98:0] addW_6600;
wire [7:0] slice_2693;
wire [45:0] concat_7356;
wire [25:0] lsl_3449;
wire [64:0] slice_4205;
wire [99:0] addW_298;
wire [15:0] mul_4961;
wire [15:0] slice_1054;
wire [15:0] mul_5717;
wire [17:0] slice_1810;
wire [15:0] slice_6473;
wire [19:0] addW_2566;
wire [66:0] concat_7229;
wire [8:0] slice_3322;
wire [195:0] concat_4078;
wire [15:0] slice_171;
wire [70:0] subW_4834;
wire [15:0] mulnw_927;
wire [39:0] mul_5590;
wire [196:0] addW_1683;
wire [15:0] slice_6346;
wire [7:0] slice_2439;
wire [31:0] slice_7102;
wire [17:0] slice_3195;
wire [31:0] slice_3951;
wire [19:0] addW_44;
wire [17:0] slice_4707;
wire [15:0] slice_800;
wire [41:0] subW_5463;
wire [7:0] slice_1556;
wire [16:0] mulnw_6219;
wire [65:0] concat_2312;
wire [17:0] add_6975;
wire [17:0] slice_3068;
wire [49:0] concat_3824;
wire [17:0] slice_4580;
wire [19:0] addW_673;
wire [133:0] concat_5336;
wire [16:0] mulnw_1429;
wire [15:0] mulnw_6092;
wire [32:0] lsl_2185;
wire [40:0] subW_6848;
wire [31:0] slice_2941;
wire [7:0] slice_3697;
wire [50:0] addW_4453;
wire [31:0] mul_546;
wire [32:0] lsl_5209;
wire [68:0] subW_1302;
wire [33:0] add_5965;
wire [15:0] mul_2058;
wire [516:0] concat_6721;
wire [63:0] slice_2814;
wire [66:0] addW_7477;
wire [25:0] lsl_3570;
wire [97:0] concat_4326;
wire [17:0] slice_419;
wire [33:0] add_5082;
wire [97:0] concat_1175;
wire [7:0] slice_5838;
wire [17:0] add_1931;
wire [34:0] addW_6594;
wire [15:0] slice_2687;
wire [13:0] slice_7350;
wire [32:0] lsl_3443;
wire [128:0] slice_4199;
wire [41:0] subW_292;
wire [7:0] slice_4955;
wire [32:0] slice_1048;
wire [7:0] slice_5711;
wire [31:0] slice_1804;
wire [25:0] lsl_6467;
wire [27:0] mul_2560;
wire [15:0] mul_7223;
wire [17:0] add_3316;
wire [67:0] subW_4072;
wire [33:0] addW_165;
wire [39:0] mul_4828;
wire [49:0] concat_921;
wire [17:0] slice_5584;
wire [71:0] subW_1677;
wire [32:0] slice_6340;
wire [15:0] slice_2433;
wire [70:0] subW_7096;
wire [31:0] slice_3189;
wire [34:0] addW_3945;
wire [35:0] mul_38;
wire [66:0] concat_4701;
wire [32:0] slice_794;
wire [17:0] slice_5457;
wire [7:0] slice_1550;
wire [15:0] slice_6213;
wire [19:0] addW_2306;
wire [16:0] mulnw_6969;
wire [19:0] addW_3062;
wire [16:0] slice_3818;
wire [31:0] slice_4574;
wire [27:0] mul_667;
wire [17:0] slice_5330;
wire [25:0] lsl_1423;
wire [49:0] concat_6086;
wire [15:0] mul_2179;
wire [35:0] mul_6842;
wire [39:0] mul_2935;
wire [1030:0] concat_7598;
wire [8:0] slice_3691;
wire [17:0] add_4447;
wire [31:0] slice_540;
wire [15:0] mul_5203;
wire [33:0] add_1296;
wire [7:0] slice_5959;
wire [7:0] slice_2052;
wire [63:0] slice_6715;
wire [99:0] addW_2808;
wire [71:0] subW_7471;
wire [32:0] lsl_3564;
wire [40:0] subW_4320;
wire [31:0] slice_413;
wire [7:0] slice_5076;
wire [40:0] subW_1169;
wire [15:0] slice_5832;
wire [16:0] mulnw_1925;
wire [15:0] mulnw_6588;
wire [33:0] addW_2681;
wire [50:0] addW_7344;
wire [15:0] mul_3437;
wire [388:0] addW_4193;
wire [17:0] slice_286;
wire [26:0] add_4949;
wire [63:0] slice_1042;
wire [15:0] slice_5705;
wire [39:0] mul_1798;
wire [32:0] lsl_6461;
wire [511:0] slice_2554;
wire [7:0] slice_7217;
wire [16:0] mulnw_3310;
wire [26:0] add_4066;
wire [41:0] subW_159;
wire [17:0] slice_4822;
wire [16:0] slice_915;
wire [34:0] addW_5578;
wire [40:0] subW_1671;
wire [98:0] addW_6334;
wire [32:0] slice_2427;
wire [39:0] mul_7090;
wire [39:0] mul_3183;
wire [15:0] mulnw_3939;
wire [13:0] slice_32;
wire [15:0] mul_4695;
wire [34:0] addW_788;
wire [31:0] slice_5451;
wire [16:0] mulnw_1544;
wire [33:0] addW_6207;
wire [17:0] slice_2300;
wire [25:0] lsl_6963;
wire [31:0] mul_3056;
wire [194:0] concat_3812;
wire [67:0] subW_4568;
wire [63:0] slice_661;
wire [19:0] addW_5324;
wire [32:0] lsl_1417;
wire [16:0] slice_6080;
wire [7:0] slice_2173;
wire [13:0] slice_6836;
wire [17:0] slice_2929;
wire [128:0] slice_7592;
wire [33:0] mul_3685;
wire [16:0] mulnw_4441;
wire [39:0] mul_534;
wire [7:0] slice_5197;
wire [7:0] slice_1290;
wire [8:0] slice_5953;
wire [26:0] add_2046;
wire [100:0] addW_6709;
wire [41:0] subW_2802;
wire [40:0] subW_7465;
wire [31:0] mul_3558;
wire [35:0] mul_4314;
wire [39:0] mul_407;
wire [8:0] slice_5070;
wire [35:0] mul_1163;
wire [32:0] slice_5826;
wire [15:0] slice_1919;
wire [8:0] slice_6582;
wire [17:0] slice_2675;
wire [17:0] add_7338;
wire [7:0] slice_3431;
wire [135:0] subW_4187;
wire [34:0] addW_280;
wire [15:0] mulnw_4943;
wire [66:0] concat_1036;
wire [32:0] slice_5699;
wire [17:0] slice_1792;
wire [15:0] mul_6455;
wire [511:0] slice_2548;
wire [26:0] add_7211;
wire [15:0] slice_3304;
wire [16:0] mulnw_4060;
wire [17:0] slice_153;
wire [34:0] addW_4816;
wire [65:0] concat_909;
wire [41:0] subW_5572;
wire [35:0] mul_1665;
wire [34:0] addW_6328;
wire [31:0] slice_2421;
wire [17:0] slice_7084;
wire [17:0] slice_3177;
wire [8:0] slice_3933;
wire [7:0] slice_4689;
wire [15:0] mulnw_782;
wire [41:0] subW_5445;
wire [7:0] slice_1538;
wire [41:0] subW_6201;
wire [66:0] concat_2294;
wire [32:0] lsl_6957;
wire [31:0] slice_3050;
wire [67:0] subW_3806;
wire [26:0] add_4562;
wire [69:0] concat_655;
wire [31:0] mul_5318;
wire [31:0] mul_1411;
wire [194:0] concat_6074;
wire [15:0] slice_2167;
wire [40:0] subW_6830;
wire [31:0] slice_2923;
wire [197:0] addW_7586;
wire [31:0] slice_3679;
wire [25:0] lsl_4435;
wire [17:0] slice_528;
wire [15:0] slice_5191;
wire [7:0] slice_1284;
wire [33:0] mul_5947;
wire [15:0] mulnw_2040;
wire [41:0] subW_6703;
wire [17:0] slice_2796;
wire [35:0] mul_7459;
wire [65:0] addW_3552;
wire [13:0] slice_4308;
wire [17:0] slice_401;
wire [33:0] mul_5064;
wire [13:0] slice_1157;
wire [34:0] addW_5820;
wire [32:0] slice_1913;
wire [17:0] add_6576;
wire [19:0] addW_2669;
wire [16:0] mulnw_7332;
wire [15:0] slice_3425;
wire [70:0] subW_4181;
wire [31:0] slice_274;
wire [49:0] concat_4937;
wire [15:0] mul_1030;
wire [31:0] slice_5693;
wire [13:0] slice_1786;
wire [7:0] slice_6449;
wire [517:0] concat_2542;
wire [15:0] mulnw_7205;
wire [32:0] slice_3298;
wire [33:0] add_4054;
wire [31:0] slice_147;
wire [41:0] subW_4810;
wire [19:0] addW_903;
wire [17:0] slice_5566;
wire [15:0] slice_1659;
wire [15:0] mulnw_6322;
wire [51:0] addW_2415;
wire [34:0] addW_7078;
wire [13:0] slice_3171;
wire [17:0] add_3927;
wire [26:0] add_4683;
wire [8:0] slice_776;
wire [17:0] slice_5439;
wire [15:0] slice_1532;
wire [17:0] slice_6195;
wire [15:0] mul_2288;
wire [31:0] mul_6951;
wire [39:0] mul_3044;
wire [26:0] add_3800;
wire [16:0] mulnw_4556;
wire [19:0] addW_649;
wire [32:0] slice_5312;
wire [64:0] slice_1405;
wire [67:0] subW_6068;
wire [32:0] slice_2161;
wire [35:0] mul_6824;
wire [39:0] mul_2917;
wire [71:0] subW_7580;
wire [39:0] mul_3673;
wire [32:0] lsl_4429;
wire [31:0] slice_522;
wire [33:0] addW_5185;
wire [16:0] mulnw_1278;
wire [31:0] slice_5941;
wire [49:0] concat_2034;
wire [17:0] slice_6697;
wire [34:0] addW_2790;
wire [15:0] slice_7453;
wire [130:0] concat_3546;
wire [40:0] subW_4302;
wire [13:0] slice_395;
wire [513:0] addW_5058;
wire [40:0] subW_1151;
wire [15:0] mulnw_5814;
wire [26:0] add_1907;
wire [16:0] mulnw_6570;
wire [27:0] mul_2663;
wire [25:0] lsl_7326;
wire [33:0] addW_3419;
wire [39:0] mul_4175;
wire [39:0] mul_268;
wire [16:0] slice_4931;
wire [7:0] slice_1024;
wire [51:0] addW_5687;
wire [71:0] subW_1780;
wire [15:0] slice_6443;
wire [64:0] slice_2536;
wire [49:0] concat_7199;
wire [26:0] add_3292;
wire [7:0] slice_4048;
wire [41:0] subW_141;
wire [17:0] slice_4804;
wire [17:0] slice_897;
wire [31:0] slice_5560;
wire [50:0] addW_1653;
wire [8:0] slice_6316;
wire [49:0] concat_2409;
wire [41:0] subW_7072;
wire [71:0] subW_3165;
wire [16:0] mulnw_3921;
wire [15:0] mulnw_4677;
wire [17:0] add_770;
wire [31:0] slice_5433;
wire [97:0] concat_1526;
wire [31:0] slice_6189;
wire [7:0] slice_2282;
wire [16:0] slice_6945;
wire [17:0] slice_3038;
wire [16:0] mulnw_3794;
wire [33:0] add_4550;
wire [17:0] slice_643;
wire [26:0] add_5306;
wire [387:0] concat_1399;
wire [26:0] add_6062;
wire [63:0] slice_2155;
wire [63:0] slice_6818;
wire [17:0] slice_2911;
wire [40:0] subW_7574;
wire [17:0] slice_3667;
wire [31:0] mul_4423;
wire [26:0] add_516;
wire [17:0] slice_5179;
wire [7:0] slice_1272;
wire [39:0] mul_5935;
wire [16:0] slice_2028;
wire [34:0] addW_6691;
wire [17:0] slice_2784;
wire [47:0] addW_7447;
wire [15:0] slice_3540;
wire [35:0] mul_4296;
wire [68:0] subW_389;
wire [513:0] addW_5052;
wire [35:0] mul_1145;
wire [8:0] slice_5808;
wire [16:0] mulnw_1901;
wire [15:0] slice_6564;
wire [17:0] slice_2657;
wire [32:0] lsl_7320;
wire [17:0] slice_3413;
wire [17:0] slice_4169;
wire [17:0] slice_262;
wire [196:0] concat_4925;
wire [26:0] add_1018;
wire [49:0] concat_5681;
wire [40:0] subW_1774;
wire [32:0] slice_6437;
wire [100:0] addW_2530;
wire [16:0] slice_7193;
wire [16:0] mulnw_3286;
wire [8:0] slice_4042;
wire [17:0] slice_135;
wire [31:0] slice_4798;
wire [65:0] concat_891;
wire [34:0] addW_5554;
wire [17:0] add_1647;
wire [17:0] add_6310;
wire [15:0] slice_2403;
wire [17:0] slice_7066;
wire [40:0] subW_3159;
wire [15:0] slice_3915;
wire [49:0] concat_4671;
wire [16:0] mulnw_764;
wire [31:0] slice_5427;
wire [40:0] subW_1520;
wire [41:0] subW_6183;
wire [26:0] add_2276;
wire [33:0] add_6939;
wire [31:0] slice_3032;
wire [33:0] add_3788;
wire [7:0] slice_4544;
wire [98:0] concat_637;
wire [16:0] mulnw_5300;
wire [132:0] subW_1393;
wire [16:0] mulnw_6056;
wire [66:0] concat_2149;
wire [99:0] addW_6812;
wire [13:0] slice_2905;
wire [35:0] mul_7568;
wire [31:0] slice_3661;
wire [16:0] slice_4417;
wire [16:0] mulnw_510;
wire [19:0] addW_5173;
wire [15:0] slice_1266;
wire [17:0] slice_5929;
wire [65:0] concat_2022;
wire [15:0] slice_6685;
wire [19:0] addW_2778;
wire [45:0] concat_7441;
wire [25:0] lsl_3534;
wire [63:0] slice_4290;
wire [33:0] add_383;
wire [255:0] slice_5046;
wire [63:0] slice_1139;
wire [17:0] add_5802;
wire [33:0] add_1895;
wire [33:0] addW_6558;
wire [19:0] addW_2651;
wire [31:0] mul_7314;
wire [19:0] addW_3407;
wire [34:0] addW_4163;
wire [31:0] slice_256;
wire [70:0] subW_4919;
wire [15:0] mulnw_1012;
wire [15:0] slice_5675;
wire [35:0] mul_1768;
wire [129:0] addW_6431;
wire [41:0] subW_2524;
wire [195:0] concat_7187;
wire [33:0] add_3280;
wire [33:0] mul_4036;
wire [31:0] slice_129;
wire [34:0] addW_4792;
wire [19:0] addW_885;
wire [15:0] mulnw_5548;
wire [16:0] mulnw_1641;
wire [16:0] mulnw_6304;
wire [65:0] concat_2397;
wire [31:0] slice_7060;
wire [35:0] mul_3153;
wire [129:0] addW_3909;
wire [16:0] slice_4665;
wire [15:0] slice_758;
wire [50:0] addW_5421;
wire [35:0] mul_1514;
wire [17:0] slice_6177;
wire [15:0] mulnw_2270;
wire [7:0] slice_6933;
wire [26:0] add_3026;
wire [7:0] slice_3782;
wire [8:0] slice_4538;
wire [40:0] subW_631;
wire [33:0] add_5294;
wire [69:0] concat_1387;
wire [33:0] add_6050;
wire [15:0] mul_2143;
wire [41:0] subW_6806;
wire [68:0] subW_2899;
wire [15:0] slice_7562;
wire [39:0] mul_3655;
wire [33:0] add_4411;
wire [33:0] add_504;
wire [27:0] mul_5167;
wire [97:0] concat_1260;
wire [31:0] slice_5923;
wire [19:0] addW_2016;
wire [25:0] lsl_6679;
wire [27:0] mul_2772;
wire [13:0] slice_7435;
wire [32:0] lsl_3528;
wire [99:0] addW_4284;
wire [7:0] slice_377;
wire [389:0] addW_5040;
wire [259:0] concat_1133;
wire [16:0] mulnw_5796;
wire [7:0] slice_1889;
wire [41:0] subW_6552;
wire [27:0] mul_2645;
wire [64:0] slice_7308;
wire [27:0] mul_3401;
wire [34:0] addW_4157;
wire [26:0] add_250;
wire [39:0] mul_4913;
wire [49:0] concat_1006;
wire [65:0] concat_5669;
wire [15:0] slice_1762;
wire [133:0] subW_6425;
wire [17:0] slice_2518;
wire [67:0] subW_7181;
wire [7:0] slice_3274;
wire [31:0] slice_4030;
wire [31:0] slice_123;
wire [15:0] mulnw_4786;
wire [17:0] slice_879;
wire [8:0] slice_5542;
wire [25:0] lsl_1635;
wire [15:0] slice_6298;
wire [19:0] addW_2391;
wire [34:0] addW_7054;
wire [15:0] slice_3147;
wire [127:0] slice_3903;
wire [194:0] concat_4659;
wire [16:0] slice_752;
wire [17:0] add_5415;
wire [13:0] slice_1508;
wire [31:0] slice_6171;
wire [49:0] concat_2264;
wire [7:0] slice_6927;
wire [16:0] mulnw_3020;
wire [8:0] slice_3776;
wire [33:0] mul_4532;
wire [35:0] mul_625;
wire [7:0] slice_5288;
wire [19:0] addW_1381;
wire [7:0] slice_6044;
wire [7:0] slice_2137;
wire [17:0] slice_6800;
wire [33:0] add_2893;
wire [50:0] addW_7556;
wire [17:0] slice_3649;
wire [7:0] slice_4405;
wire [7:0] slice_498;
wire [17:0] slice_5161;
wire [40:0] subW_1254;
wire [39:0] mul_5917;
wire [17:0] slice_2010;
wire [32:0] lsl_6673;
wire [15:0] slice_2766;
wire [50:0] addW_7429;
wire [15:0] mul_3522;
wire [41:0] subW_4278;
wire [7:0] slice_371;
wire [135:0] subW_5034;
wire [31:0] slice_1127;
wire [15:0] slice_5790;
wire [8:0] slice_1883;
wire [17:0] slice_6546;
wire [63:0] slice_2639;
wire [17:0] slice_3395;
wire [15:0] mulnw_4151;
wire [16:0] mulnw_244;
wire [17:0] slice_4907;
wire [16:0] slice_1000;
wire [19:0] addW_5663;
wire [47:0] addW_1756;
wire [70:0] subW_6419;
wire [34:0] addW_2512;
wire [26:0] add_7175;
wire [8:0] slice_3268;
wire [39:0] mul_4024;
wire [50:0] addW_117;
wire [8:0] slice_4780;
wire [255:0] slice_873;
wire [17:0] add_5536;
wire [32:0] lsl_1629;
wire [33:0] addW_6292;
wire [17:0] slice_2385;
wire [15:0] mulnw_7048;
wire [47:0] addW_3141;
wire [131:0] concat_3897;
wire [67:0] subW_4653;
wire [63:0] slice_746;
wire [16:0] mulnw_5409;
wire [40:0] subW_1502;
wire [127:0] slice_6165;
wire [16:0] slice_2258;
wire [16:0] mulnw_6921;
wire [33:0] add_3014;
wire [33:0] mul_3770;
wire [31:0] slice_4526;
wire [13:0] slice_619;
wire [8:0] slice_5282;
wire [17:0] slice_1375;
wire [8:0] slice_6038;
wire [26:0] add_2131;
wire [34:0] addW_6794;
wire [7:0] slice_2887;
wire [17:0] add_7550;
wire [127:0] slice_3643;
wire [7:0] slice_4399;
wire [8:0] slice_492;
wire [19:0] addW_5155;
wire [35:0] mul_1248;
wire [17:0] slice_5911;
wire [65:0] concat_2004;
wire [15:0] mul_6667;
wire [25:0] lsl_2760;
wire [17:0] add_7423;
wire [7:0] slice_3516;
wire [17:0] slice_4272;
wire [16:0] mulnw_365;
wire [70:0] subW_5028;
wire [51:0] addW_1121;
wire [16:0] slice_5784;
wire [33:0] mul_1877;
wire [31:0] slice_6540;
wire [66:0] concat_2633;
wire [135:0] subW_7296;
wire [19:0] addW_3389;
wire [8:0] slice_4145;
wire [33:0] add_238;
wire [34:0] addW_4901;
wire [65:0] concat_994;
wire [17:0] slice_5657;
wire [45:0] concat_1750;
wire [39:0] mul_6413;
wire [15:0] slice_2506;
wire [16:0] mulnw_7169;
wire [33:0] mul_3262;
wire [17:0] slice_4018;
wire [17:0] add_111;
wire [17:0] add_4774;
wire [516:0] concat_867;
wire [16:0] mulnw_5530;
wire [31:0] mul_1623;
wire [41:0] subW_6286;
wire [66:0] concat_2379;
wire [8:0] slice_7042;
wire [45:0] concat_3135;
wire [17:0] slice_3891;
wire [26:0] add_4647;
wire [66:0] concat_740;
wire [25:0] lsl_5403;
wire [35:0] mul_1496;
wire [131:0] concat_6159;
wire [64:0] slice_2252;
wire [7:0] slice_6915;
wire [7:0] slice_3008;
wire [31:0] slice_3764;
wire [39:0] mul_4520;
wire [33:0] add_613;
wire [33:0] mul_5276;
wire [98:0] concat_1369;
wire [33:0] mul_6032;
wire [15:0] mulnw_2125;
wire [17:0] slice_6788;
wire [7:0] slice_2881;
wire [16:0] mulnw_7544;
wire [63:0] slice_3637;
wire [16:0] mulnw_4393;
wire [33:0] mul_486;
wire [27:0] mul_5149;
wire [13:0] slice_1242;
wire [127:0] slice_5905;
wire [19:0] addW_1998;
wire [7:0] slice_6661;
wire [32:0] lsl_2754;
wire [16:0] mulnw_7417;
wire [15:0] slice_3510;
wire [34:0] addW_4266;
wire [7:0] slice_359;
wire [39:0] mul_5022;
wire [49:0] concat_1115;
wire [31:0] slice_5778;
wire [66:0] addW_1871;
wire [41:0] subW_6534;
wire [15:0] mul_2627;
wire [70:0] subW_7290;
wire [27:0] mul_3383;
wire [17:0] add_4139;
wire [7:0] slice_232;
wire [41:0] subW_4895;
wire [19:0] addW_988;
wire [66:0] concat_5651;
wire [13:0] slice_1744;
wire [17:0] slice_6407;
wire [25:0] lsl_2500;
wire [33:0] add_7163;
wire [66:0] addW_3256;
wire [31:0] slice_4012;
wire [16:0] mulnw_105;
wire [16:0] mulnw_4768;
wire [63:0] slice_861;
wire [15:0] slice_5524;
wire [16:0] slice_1617;
wire [17:0] slice_6280;
wire [15:0] mul_2373;
wire [17:0] add_7036;
wire [13:0] slice_3129;
wire [19:0] addW_3885;
wire [16:0] mulnw_4641;
wire [15:0] mul_734;
wire [32:0] lsl_5397;
wire [63:0] slice_1490;
wire [17:0] slice_6153;
wire [259:0] concat_2246;
wire [15:0] slice_6909;
wire [8:0] slice_3002;
wire [39:0] mul_3758;
wire [17:0] slice_4514;
wire [7:0] slice_607;
wire [15:0] slice_5270;
wire [40:0] subW_1363;
wire [31:0] slice_6026;
wire [49:0] concat_2119;
wire [19:0] addW_6782;
wire [16:0] mulnw_2875;
wire [25:0] lsl_7538;
wire [99:0] addW_3631;
wire [7:0] slice_4387;
wire [65:0] addW_480;
wire [63:0] slice_5143;
wire [40:0] subW_1236;
wire [255:0] slice_5899;
wire [17:0] slice_1992;
wire [15:0] slice_6655;
wire [15:0] mul_2748;
wire [25:0] lsl_7411;
wire [33:0] addW_3504;
wire [17:0] slice_4260;
wire [15:0] slice_353;
wire [17:0] slice_5016;
wire [15:0] slice_1109;
wire [51:0] addW_5772;
wire [68:0] subW_1865;
wire [17:0] slice_6528;
wire [7:0] slice_2621;
wire [39:0] mul_7284;
wire [13:0] slice_3377;
wire [16:0] mulnw_4133;
wire [8:0] slice_226;
wire [17:0] slice_4889;
wire [17:0] slice_982;
wire [15:0] mul_5645;
wire [50:0] addW_1738;
wire [34:0] addW_6401;
wire [32:0] lsl_2494;
wire [7:0] slice_7157;
wire [68:0] subW_3250;
wire [39:0] mul_4006;
wire [25:0] lsl_99;
wire [15:0] slice_4762;
wire [100:0] addW_855;
wire [16:0] slice_5518;
wire [33:0] add_1611;
wire [31:0] slice_6274;
wire [7:0] slice_2367;
wire [16:0] mulnw_7030;
wire [50:0] addW_3123;
wire [31:0] mul_3879;
wire [33:0] add_4635;
wire [7:0] slice_728;
wire [31:0] mul_5391;
wire [99:0] addW_1484;
wire [19:0] addW_6147;
wire [31:0] slice_2240;
wire [32:0] slice_6903;
wire [33:0] mul_2996;
wire [17:0] slice_3752;
wire [31:0] slice_4508;
wire [7:0] slice_601;
wire [25:0] lsl_5264;
wire [35:0] mul_1357;
wire [39:0] mul_6020;
wire [16:0] slice_2113;
wire [27:0] mul_6776;
wire [7:0] slice_2869;
wire [32:0] lsl_7532;
wire [41:0] subW_3625;
wire [15:0] slice_4381;
wire [68:0] subW_474;
wire [69:0] concat_5137;
wire [35:0] mul_1230;
wire [262:0] concat_5893;
wire [13:0] slice_1986;
wire [32:0] slice_6649;
wire [7:0] slice_2742;
wire [32:0] lsl_7405;
wire [17:0] slice_3498;
wire [19:0] addW_4254;
wire [97:0] concat_347;
wire [34:0] addW_5010;
wire [65:0] concat_1103;
wire [49:0] concat_5766;
wire [33:0] add_1859;
wire [31:0] slice_6522;
wire [26:0] add_2615;
wire [17:0] slice_7278;
wire [127:0] slice_3371;
wire [15:0] slice_4127;
wire [33:0] mul_220;
wire [31:0] slice_4883;
wire [65:0] concat_976;
wire [7:0] slice_5639;
wire [17:0] add_1732;
wire [41:0] subW_6395;
wire [15:0] mul_2488;
wire [8:0] slice_7151;
wire [33:0] add_3244;
wire [17:0] slice_4000;
wire [130:0] addW_4756;
wire [41:0] subW_849;
wire [31:0] slice_5512;
wire [7:0] slice_1605;
wire [41:0] subW_6268;
wire [26:0] add_2361;
wire [15:0] slice_7024;
wire [17:0] add_3117;
wire [31:0] slice_3873;
wire [7:0] slice_4629;
wire [26:0] add_722;
wire [16:0] slice_5385;
wire [41:0] subW_1478;
wire [31:0] mul_6141;
wire [51:0] addW_2234;
wire [98:0] addW_6897;
wire [65:0] addW_2990;
wire [31:0] slice_3746;
wire [39:0] mul_4502;
wire [16:0] mulnw_595;
wire [32:0] lsl_5258;
wire [13:0] slice_1351;
wire [17:0] slice_6014;
wire [65:0] concat_2107;
wire [15:0] slice_6770;
wire [15:0] slice_2863;
wire [31:0] mul_7526;
wire [17:0] slice_3619;
wire [32:0] slice_4375;
wire [33:0] add_468;
wire [19:0] addW_5131;
wire [63:0] slice_1224;
wire [32:0] slice_5887;
wire [196:0] addW_1980;
wire [34:0] addW_6643;
wire [15:0] slice_2736;
wire [31:0] mul_7399;
wire [19:0] addW_3492;
wire [27:0] mul_4248;
wire [40:0] subW_341;
wire [34:0] addW_5004;
wire [19:0] addW_1097;
wire [15:0] slice_5760;
wire [7:0] slice_1853;
wire [31:0] slice_6516;
wire [15:0] mulnw_2609;
wire [34:0] addW_7272;
wire [196:0] addW_3365;
wire [32:0] slice_4121;
wire [65:0] addW_214;
wire [34:0] addW_4877;
wire [19:0] addW_970;
wire [26:0] add_5633;
wire [16:0] mulnw_1726;
wire [17:0] slice_6389;
wire [7:0] slice_2482;
wire [33:0] mul_7145;
wire [7:0] slice_3238;
wire [13:0] slice_3994;
wire [127:0] slice_4750;
wire [17:0] slice_843;
wire [50:0] addW_5506;
wire [7:0] slice_1599;
wire [17:0] slice_6262;
wire [15:0] mulnw_2355;
wire [128:0] slice_7018;
wire [16:0] mulnw_3111;
wire [39:0] mul_3867;
wire [8:0] slice_4623;
wire [15:0] mulnw_716;
wire [47:0] addW_5379;
wire [17:0] slice_1472;
wire [31:0] slice_6135;
wire [49:0] concat_2228;
wire [34:0] addW_6891;
wire [68:0] subW_2984;
wire [39:0] mul_3740;
wire [17:0] slice_4496;
wire [7:0] slice_589;
wire [15:0] mul_5252;
wire [33:0] add_1345;
wire [31:0] slice_6008;
wire [19:0] addW_2101;
wire [25:0] lsl_6764;
wire [97:0] concat_2857;
wire [16:0] slice_7520;
wire [34:0] addW_3613;
wire [98:0] addW_4369;
wire [7:0] slice_462;
wire [17:0] slice_5125;
wire [98:0] addW_1218;
wire [51:0] addW_5881;
wire [71:0] subW_1974;
wire [15:0] mulnw_6637;
wire [32:0] slice_2730;
wire [64:0] slice_7393;
wire [27:0] mul_3486;
wire [15:0] slice_4242;
wire [35:0] mul_335;
wire [15:0] mulnw_4998;
wire [17:0] slice_1091;
wire [65:0] concat_5754;
wire [7:0] slice_1847;
wire [51:0] addW_6510;
wire [49:0] concat_2603;
wire [34:0] addW_7266;
wire [71:0] subW_3359;
wire [26:0] add_4115;
wire [31:0] slice_208;
wire [15:0] mulnw_4871;
wire [17:0] slice_964;
wire [15:0] mulnw_5627;
wire [25:0] lsl_1720;
wire [31:0] slice_6383;
wire [15:0] slice_2476;
wire [31:0] slice_7139;
wire [7:0] slice_3232;
wire [71:0] subW_3988;
wire [131:0] concat_4744;
wire [34:0] addW_837;
wire [17:0] add_5500;
wire [16:0] mulnw_1593;
wire [31:0] slice_6256;
wire [49:0] concat_2349;
wire [63:0] slice_7012;
wire [25:0] lsl_3105;
wire [17:0] slice_3861;
wire [33:0] mul_4617;
wire [49:0] concat_710;
wire [45:0] concat_5373;
wire [34:0] addW_1466;
wire [39:0] mul_6129;
wire [15:0] slice_2222;
wire [15:0] mulnw_6885;
wire [33:0] add_2978;
wire [17:0] slice_3734;
wire [127:0] slice_4490;
wire [15:0] slice_583;
wire [7:0] slice_5246;
wire [7:0] slice_1339;
wire [39:0] mul_6002;
wire [17:0] slice_2095;
wire [32:0] lsl_6758;
wire [40:0] subW_2851;
wire [33:0] add_7514;
wire [17:0] slice_3607;
wire [34:0] addW_4363;
wire [7:0] slice_456;
wire [98:0] concat_5119;
wire [34:0] addW_1212;
wire [49:0] concat_5875;
wire [40:0] subW_1968;
wire [8:0] slice_6631;
wire [63:0] slice_2724;
wire [99:0] addW_7387;
wire [17:0] slice_3480;
wire [25:0] lsl_4236;
wire [13:0] slice_329;
wire [8:0] slice_4992;
wire [66:0] concat_1085;
wire [19:0] addW_5748;
wire [16:0] mulnw_1841;
wire [49:0] concat_6504;
wire [16:0] slice_2597;
wire [15:0] mulnw_7260;
wire [40:0] subW_3353;
wire [16:0] mulnw_4109;
wire [50:0] addW_202;
wire [8:0] slice_4865;
wire [31:0] slice_958;
wire [49:0] concat_5621;
wire [32:0] lsl_1714;
wire [34:0] addW_6377;
wire [32:0] slice_2470;
wire [39:0] mul_7133;
wire [16:0] mulnw_3226;
wire [40:0] subW_3982;
wire [33:0] addW_75;
wire [17:0] slice_4738;
wire [66:0] concat_831;
wire [16:0] mulnw_5494;
wire [7:0] slice_1587;
wire [31:0] slice_6250;
wire [16:0] slice_2343;
wire [100:0] addW_7006;
wire [32:0] lsl_3099;
wire [31:0] slice_3855;
wire [31:0] slice_4611;
wire [16:0] slice_704;
wire [13:0] slice_5367;
wire [17:0] slice_1460;
wire [17:0] slice_6123;
wire [65:0] concat_2216;
wire [8:0] slice_6879;
wire [7:0] slice_2972;
wire [13:0] slice_3728;
wire [63:0] slice_4484;
wire [16:0] slice_577;
wire [15:0] slice_5240;
wire [7:0] slice_1333;
wire [17:0] slice_5996;
wire [65:0] concat_2089;
wire [15:0] mul_6752;
wire [35:0] mul_2845;
wire [7:0] slice_7508;
wire [19:0] addW_3601;
wire [15:0] mulnw_4357;
wire [16:0] mulnw_450;
wire [40:0] subW_5113;
wire [15:0] mulnw_1206;
wire [15:0] slice_5869;
wire [35:0] mul_1962;
wire [17:0] add_6625;
wire [66:0] concat_2718;
wire [41:0] subW_7381;
wire [19:0] addW_3474;
wire [32:0] lsl_4230;
wire [40:0] subW_323;
wire [17:0] add_4986;
wire [15:0] mul_1079;
wire [17:0] slice_5742;
wire [7:0] slice_1835;
wire [15:0] slice_6498;
wire [65:0] concat_2591;
wire [8:0] slice_7254;
wire [35:0] mul_3347;
wire [33:0] add_4103;
wire [17:0] add_196;
wire [17:0] add_4859;
wire [67:0] subW_952;
wire [16:0] slice_5615;
wire [31:0] mul_1708;
wire [15:0] mulnw_6371;
wire [34:0] addW_2464;
wire [17:0] slice_7127;
wire [7:0] slice_3220;
wire [35:0] mul_3976;
wire [65:0] concat_69;
wire [19:0] addW_4732;
wire [15:0] mul_825;
wire [25:0] lsl_5488;
wire [15:0] slice_1581;
wire [50:0] addW_6244;
wire [131:0] concat_2337;
wire [41:0] subW_7000;
wire [31:0] mul_3093;
wire [26:0] add_3849;
wire [39:0] mul_4605;
wire [65:0] concat_698;
wire [47:0] addW_5361;
wire [19:0] addW_1454;
wire [31:0] slice_6117;
wire [19:0] addW_2210;
wire [17:0] add_6873;
wire [7:0] slice_2966;
wire [68:0] subW_3722;
wire [100:0] addW_4478;
wire [387:0] concat_571;
wire [32:0] slice_5234;
wire [16:0] mulnw_1327;
wire [13:0] slice_5990;
wire [19:0] addW_2083;
wire [7:0] slice_6746;
wire [13:0] slice_2839;
wire [7:0] slice_7502;
wire [27:0] mul_3595;
wire [8:0] slice_4351;
wire [7:0] slice_444;
wire [35:0] mul_5107;
wire [8:0] slice_1200;
wire [66:0] concat_5863;
wire [15:0] slice_1956;
wire [16:0] mulnw_6619;
wire [15:0] mul_2712;
wire [17:0] slice_7375;
wire [27:0] mul_3468;
wire [15:0] mul_4224;
wire [35:0] mul_317;
wire [16:0] mulnw_4980;
wire [7:0] slice_1073;
wire [66:0] concat_5736;
wire [15:0] slice_1829;
wire [65:0] concat_6492;
wire [19:0] addW_2585;
wire [17:0] add_7248;
wire [15:0] slice_3341;
wire [7:0] slice_4097;
wire [16:0] mulnw_190;
wire [16:0] mulnw_4853;
wire [26:0] add_946;
wire [64:0] slice_5609;
wire [64:0] slice_1702;
wire [8:0] slice_6365;
wire [15:0] mulnw_2458;
wire [31:0] slice_7121;
wire [15:0] slice_3214;
wire [15:0] slice_3970;
wire [19:0] addW_63;
wire [31:0] mul_4726;
wire [7:0] slice_819;
wire [32:0] lsl_5482;
wire [32:0] slice_1575;
wire [17:0] add_6238;
wire [17:0] slice_2331;
wire [17:0] slice_6994;
wire [64:0] slice_3087;
wire [16:0] mulnw_3843;
wire [17:0] slice_4599;
wire [19:0] addW_692;
wire [45:0] concat_5355;
wire [27:0] mul_1448;
wire [26:0] add_6111;
wire [17:0] slice_2204;
wire [16:0] mulnw_6867;
wire [16:0] mulnw_2960;
wire [33:0] add_3716;
wire [41:0] subW_4472;
wire [132:0] subW_565;
wire [63:0] slice_5228;
wire [7:0] slice_1321;
wire [68:0] subW_5984;
wire [17:0] slice_2077;
wire [15:0] slice_6740;
wire [40:0] subW_2833;
wire [16:0] mulnw_7496;
wire [15:0] slice_3589;
wire [17:0] add_4345;
wire [15:0] slice_438;
wire [13:0] slice_5101;
wire [17:0] add_1194;
wire [15:0] mul_5857;
wire [50:0] addW_1950;
wire [15:0] slice_6613;
wire [7:0] slice_2706;
wire [34:0] addW_7369;
wire [63:0] slice_3462;
wire [7:0] slice_4218;
wire [63:0] slice_311;
wire [15:0] slice_4974;
wire [26:0] add_1067;
wire [15:0] mul_5730;
wire [97:0] concat_1823;
wire [19:0] addW_6486;
wire [17:0] slice_2579;
wire [16:0] mulnw_7242;
wire [50:0] addW_3335;
wire [8:0] slice_4091;
wire [25:0] lsl_184;
wire [15:0] slice_4847;
wire [16:0] mulnw_940;
wire [195:0] addW_5603;
wire [128:0] slice_1696;
wire [17:0] add_6359;
wire [8:0] slice_2452;
wire [39:0] mul_7115;
wire [97:0] concat_3208;
wire [47:0] addW_3964;
wire [17:0] slice_57;
wire [31:0] slice_4720;
wire [26:0] add_813;
wire [31:0] mul_5476;
wire [98:0] addW_1569;
wire [16:0] mulnw_6232;
wire [19:0] addW_2325;
wire [34:0] addW_6988;
wire [387:0] concat_3081;
wire [33:0] add_3837;
wire [31:0] slice_4593;
wire [17:0] slice_686;
wire [13:0] slice_5349;
wire [15:0] slice_1442;
wire [16:0] mulnw_6105;
wire [66:0] concat_2198;
wire [15:0] slice_6861;
wire [7:0] slice_2954;
wire [7:0] slice_3710;
wire [17:0] slice_4466;
wire [69:0] concat_559;
wire [66:0] concat_5222;
wire [15:0] slice_1315;
wire [33:0] add_5978;
wire [31:0] slice_2071;
wire [32:0] slice_6734;
wire [35:0] mul_2827;
wire [7:0] slice_7490;
wire [25:0] lsl_3583;
wire [16:0] mulnw_4339;
wire [97:0] concat_432;
wire [33:0] add_5095;
wire [16:0] mulnw_1188;
wire [7:0] slice_5851;
wire [17:0] add_1944;
wire [16:0] slice_6607;
wire [26:0] add_2700;
wire [17:0] slice_7363;
wire [66:0] concat_3456;
wire [15:0] slice_4212;
wire [259:0] concat_305;
wire [32:0] slice_4968;
wire [15:0] mulnw_1061;
wire [7:0] slice_5724;
wire [40:0] subW_1817;
wire [17:0] slice_6480;
wire [65:0] concat_2573;
wire [15:0] slice_7236;
wire [17:0] add_3329;
wire [33:0] mul_4085;
wire [32:0] lsl_178;
wire [16:0] slice_4841;
wire [33:0] add_934;
wire [71:0] subW_5597;
wire [516:0] concat_1690;
wire [16:0] mulnw_6353;
wire [17:0] add_2446;
wire [17:0] slice_7109;
wire [40:0] subW_3202;
wire [45:0] concat_3958;
wire [65:0] concat_51;
wire [39:0] mul_4714;
wire [15:0] mulnw_807;
wire [16:0] slice_5470;
wire [34:0] addW_1563;
wire [25:0] lsl_6226;
wire [31:0] mul_2319;
wire [15:0] slice_6982;
wire [132:0] subW_3075;
wire [7:0] slice_3831;
wire [39:0] mul_4587;
wire [65:0] concat_680;
wire [63:0] slice_5343;
wire [25:0] lsl_1436;
wire [33:0] add_6099;
wire [15:0] mul_2192;
wire [33:0] addW_6855;
wire [15:0] slice_2948;
wire [7:0] slice_3704;
wire [34:0] addW_4460;
wire [19:0] addW_553;
wire [15:0] mul_5216;
wire [32:0] slice_1309;
wire [7:0] slice_5972;
wire [67:0] subW_2065;
wire [64:0] slice_6728;
wire [63:0] slice_2821;
wire [15:0] slice_7484;
wire [32:0] lsl_3577;
wire [15:0] slice_4333;
wire [40:0] subW_426;
wire [7:0] slice_5089;
wire [15:0] slice_1182;
wire [26:0] add_5845;
wire [16:0] mulnw_1938;
wire [31:0] slice_6601;
wire [15:0] mulnw_2694;
wire [19:0] addW_7357;
wire [15:0] mul_3450;
wire [32:0] slice_4206;
wire [31:0] slice_299;
wire [26:0] add_4962;
wire [49:0] concat_1055;
wire [26:0] add_5718;
wire [35:0] mul_1811;
wire [66:0] concat_6474;
wire [19:0] addW_2567;
wire [32:0] slice_7230;
wire [16:0] mulnw_3323;
wire [66:0] addW_4079;
wire [31:0] mul_172;
wire [71:0] subW_4835;
wire [7:0] slice_928;
wire [40:0] subW_5591;
wire [63:0] slice_1684;
wire [15:0] slice_6347;
wire [16:0] mulnw_2440;
wire [13:0] slice_7103;
wire [35:0] mul_3196;
wire [13:0] slice_3952;
wire [19:0] addW_45;
wire [17:0] slice_4708;
wire [49:0] concat_801;
wire [47:0] addW_5464;
wire [15:0] mulnw_1557;
wire [32:0] lsl_6220;
wire [31:0] slice_2313;
wire [25:0] lsl_6976;
wire [69:0] concat_3069;
wire [8:0] slice_3825;
wire [17:0] slice_4581;
wire [19:0] addW_674;
wire [134:0] subW_5337;
wire [32:0] lsl_1430;
wire [7:0] slice_6093;
wire [7:0] slice_2186;
wire [41:0] subW_6849;
wire [97:0] concat_2942;
wire [16:0] mulnw_3698;
wire [15:0] slice_4454;
wire [17:0] slice_547;
wire [7:0] slice_5210;
wire [98:0] addW_1303;
wire [7:0] slice_5966;
wire [26:0] add_2059;
wire [255:0] slice_6722;
wire [259:0] concat_2815;
wire [32:0] slice_7478;
wire [15:0] mul_3571;
wire [33:0] addW_4327;
wire [35:0] mul_420;
wire [7:0] slice_5083;
wire [33:0] addW_1176;
wire [15:0] mulnw_5839;
wire [25:0] lsl_1932;
wire [50:0] addW_6595;
wire [49:0] concat_2688;
wire [27:0] mul_7351;
wire [7:0] slice_3444;
wire [64:0] slice_4200;
wire [51:0] addW_293;
wire [16:0] mulnw_4956;
wire [16:0] slice_1049;
wire [15:0] mulnw_5712;
wire [13:0] slice_1805;
wire [15:0] mul_6468;
wire [17:0] slice_2561;
wire [26:0] add_7224;
wire [25:0] lsl_3317;
wire [68:0] subW_4073;
wire [16:0] slice_166;
wire [40:0] subW_4829;
wire [8:0] slice_922;
wire [35:0] mul_5585;
wire [100:0] addW_1678;
wire [16:0] slice_6341;
wire [15:0] slice_2434;
wire [71:0] subW_7097;
wire [13:0] slice_3190;
wire [50:0] addW_3946;
wire [31:0] slice_4702;
wire [16:0] slice_795;
wire [45:0] concat_5458;
wire [8:0] slice_1551;
wire [31:0] mul_6214;
wire [39:0] mul_2307;
wire [32:0] lsl_6970;
wire [19:0] addW_3063;
wire [33:0] mul_3819;
wire [13:0] slice_4575;
wire [17:0] slice_668;
wire [69:0] concat_5331;
wire [15:0] mul_1424;
wire [8:0] slice_6087;
wire [26:0] add_2180;
wire [17:0] slice_6843;
wire [40:0] subW_2936;
wire [1031:0] subW_7599;
wire [7:0] slice_3692;
wire [25:0] lsl_4448;
wire [98:0] concat_541;
wire [26:0] add_5204;
wire [34:0] addW_1297;
wire [16:0] mulnw_5960;
wire [16:0] mulnw_2053;
wire [260:0] concat_6716;
wire [31:0] slice_2809;
wire [99:0] addW_7472;
wire [7:0] slice_3565;
wire [41:0] subW_4321;
wire [13:0] slice_414;
wire [16:0] mulnw_5077;
wire [41:0] subW_1170;
wire [49:0] concat_5833;
wire [32:0] lsl_1926;
wire [17:0] add_6589;
wire [16:0] slice_2682;
wire [15:0] slice_7345;
wire [26:0] add_3438;
wire [127:0] slice_4194;
wire [49:0] concat_287;
wire [33:0] add_4950;
wire [194:0] concat_1043;
wire [49:0] concat_5706;
wire [40:0] subW_1799;
wire [7:0] slice_6462;
wire [255:0] slice_2555;
wire [16:0] mulnw_7218;
wire [32:0] lsl_3311;
wire [33:0] add_4067;
wire [47:0] addW_160;
wire [35:0] mul_4823;
wire [33:0] mul_916;
wire [15:0] slice_5579;
wire [41:0] subW_1672;
wire [31:0] slice_6335;
wire [16:0] slice_2428;
wire [40:0] subW_7091;
wire [40:0] subW_3184;
wire [17:0] add_3940;
wire [27:0] mul_33;
wire [26:0] add_4696;
wire [50:0] addW_789;
wire [13:0] slice_5452;
wire [17:0] add_1545;
wire [16:0] slice_6208;
wire [17:0] slice_2301;
wire [15:0] mul_6964;
wire [17:0] slice_3057;
wire [65:0] addW_3813;
wire [68:0] subW_4569;
wire [31:0] slice_662;
wire [19:0] addW_5325;
wire [7:0] slice_1418;
wire [33:0] mul_6081;
wire [15:0] mulnw_2174;
wire [31:0] slice_6837;
wire [35:0] mul_2930;
wire [519:0] concat_7593;
wire [15:0] slice_3686;
wire [32:0] lsl_4442;
wire [40:0] subW_535;
wire [15:0] mulnw_5198;
wire [15:0] mulnw_1291;
wire [7:0] slice_5954;
wire [33:0] add_2047;
wire [32:0] slice_6710;
wire [51:0] addW_2803;
wire [41:0] subW_7466;
wire [15:0] slice_3559;
wire [17:0] slice_4315;
wire [40:0] subW_408;
wire [7:0] slice_5071;
wire [17:0] slice_1164;
wire [16:0] slice_5827;
wire [31:0] mul_1920;
wire [16:0] mulnw_6583;
wire [65:0] concat_2676;
wire [25:0] lsl_7339;
wire [15:0] mulnw_3432;
wire [196:0] addW_4188;
wire [15:0] slice_281;
wire [7:0] slice_4944;
wire [67:0] subW_1037;
wire [16:0] slice_5700;
wire [35:0] mul_1793;
wire [26:0] add_6456;
wire [255:0] slice_2549;
wire [33:0] add_7212;
wire [31:0] mul_3305;
wire [7:0] slice_4061;
wire [45:0] concat_154;
wire [15:0] slice_4817;
wire [31:0] slice_910;
wire [47:0] addW_5573;
wire [17:0] slice_1666;
wire [50:0] addW_6329;
wire [131:0] concat_2422;
wire [35:0] mul_7085;
wire [35:0] mul_3178;
wire [16:0] mulnw_3934;
wire [511:0] slice_27;
wire [16:0] mulnw_4690;
wire [17:0] add_783;
wire [47:0] addW_5446;
wire [16:0] mulnw_1539;
wire [47:0] addW_6202;
wire [31:0] slice_2295;
wire [7:0] slice_6958;
wire [98:0] concat_3051;
wire [68:0] subW_3807;
wire [33:0] add_4563;
wire [70:0] subW_656;
wire [17:0] slice_5319;
wire [15:0] slice_1412;
wire [65:0] addW_6075;
wire [49:0] concat_2168;
wire [41:0] subW_6831;
wire [13:0] slice_2924;
wire [64:0] slice_7587;
wire [97:0] concat_3680;
wire [15:0] mul_4436;
wire [35:0] mul_529;
wire [49:0] concat_5192;
wire [8:0] slice_1285;
wire [15:0] slice_5948;
wire [7:0] slice_2041;
wire [51:0] addW_6704;
wire [49:0] concat_2797;
wire [17:0] slice_7460;
wire [32:0] slice_3553;
wire [31:0] slice_4309;
wire [35:0] mul_402;
wire [15:0] slice_5065;
wire [31:0] slice_1158;
wire [50:0] addW_5821;
wire [16:0] slice_1914;
wire [25:0] lsl_6577;
wire [19:0] addW_2670;
wire [32:0] lsl_7333;
wire [49:0] concat_3426;
wire [71:0] subW_4182;
wire [98:0] concat_275;
wire [8:0] slice_4938;
wire [26:0] add_1031;
wire [131:0] concat_5694;
wire [63:0] slice_1787;
wire [15:0] mulnw_6450;
wire [518:0] subW_2543;
wire [7:0] slice_7206;
wire [16:0] slice_3299;
wire [7:0] slice_4055;
wire [13:0] slice_148;
wire [47:0] addW_4811;
wire [39:0] mul_904;
wire [45:0] concat_5567;
wire [34:0] addW_1660;
wire [17:0] add_6323;
wire [17:0] slice_2416;
wire [15:0] slice_7079;
wire [63:0] slice_3172;
wire [25:0] lsl_3928;
wire [33:0] add_4684;
wire [16:0] mulnw_777;
wire [45:0] concat_5440;
wire [15:0] slice_1533;
wire [45:0] concat_6196;
wire [26:0] add_2289;
wire [15:0] slice_6952;
wire [40:0] subW_3045;
wire [33:0] add_3801;
wire [7:0] slice_4557;
wire [39:0] mul_650;
wire [99:0] concat_5313;
wire [32:0] slice_1406;
wire [68:0] subW_6069;
wire [16:0] slice_2162;
wire [17:0] slice_6825;
wire [40:0] subW_2918;
wire [100:0] addW_7581;
wire [40:0] subW_3674;
wire [7:0] slice_4430;
wire [13:0] slice_523;
wire [16:0] slice_5186;
wire [17:0] add_1279;
wire [97:0] concat_5942;
wire [8:0] slice_2035;
wire [49:0] concat_6698;
wire [15:0] slice_2791;
wire [34:0] addW_7454;
wire [63:0] slice_3547;
wire [41:0] subW_4303;
wire [63:0] slice_396;
wire [256:0] slice_5059;
wire [41:0] subW_1152;
wire [17:0] add_5815;
wire [33:0] add_1908;
wire [32:0] lsl_6571;
wire [17:0] slice_2664;
wire [15:0] mul_7327;
wire [16:0] slice_3420;
wire [40:0] subW_4176;
wire [40:0] subW_269;
wire [33:0] mul_4932;
wire [16:0] mulnw_1025;
wire [17:0] slice_5688;
wire [99:0] addW_1781;
wire [49:0] concat_6444;
wire [262:0] concat_2537;
wire [8:0] slice_7200;
wire [33:0] add_3293;
wire [16:0] mulnw_4049;
wire [47:0] addW_142;
wire [45:0] concat_4805;
wire [17:0] slice_898;
wire [13:0] slice_5561;
wire [15:0] slice_1654;
wire [16:0] mulnw_6317;
wire [19:0] addW_2410;
wire [47:0] addW_7073;
wire [99:0] addW_3166;
wire [32:0] lsl_3922;
wire [7:0] slice_4678;
wire [25:0] lsl_771;
wire [13:0] slice_5434;
wire [33:0] addW_1527;
wire [13:0] slice_6190;
wire [16:0] mulnw_2283;
wire [32:0] slice_6946;
wire [35:0] mul_3039;
wire [7:0] slice_3795;
wire [7:0] slice_4551;
wire [17:0] slice_644;
wire [33:0] add_5307;
wire [129:0] addW_1400;
wire [33:0] add_6063;
wire [194:0] concat_2156;
wire [31:0] slice_6819;
wire [35:0] mul_2912;
wire [41:0] subW_7575;
wire [35:0] mul_3668;
wire [15:0] slice_4424;
wire [33:0] add_517;
wire [65:0] concat_5180;
wire [16:0] mulnw_1273;
wire [40:0] subW_5936;
wire [33:0] mul_2029;
wire [15:0] slice_6692;
wire [65:0] concat_2785;
wire [17:0] slice_7448;
wire [66:0] concat_3541;
wire [17:0] slice_4297;
wire [98:0] addW_390;
wire [256:0] slice_5053;
wire [17:0] slice_1146;
wire [16:0] mulnw_5809;
wire [7:0] slice_1902;
wire [31:0] mul_6565;
wire [65:0] concat_2658;
wire [7:0] slice_7321;
wire [65:0] concat_3414;
wire [35:0] mul_4170;
wire [35:0] mul_263;
wire [66:0] addW_4926;
wire [33:0] add_1019;
wire [19:0] addW_5682;
wire [41:0] subW_1775;
wire [16:0] slice_6438;
wire [32:0] slice_2531;
wire [33:0] mul_7194;
wire [7:0] slice_3287;
wire [7:0] slice_4043;
wire [45:0] concat_136;
wire [13:0] slice_4799;
wire [31:0] slice_892;
wire [50:0] addW_5555;
wire [25:0] lsl_1648;
wire [25:0] lsl_6311;
wire [31:0] mul_2404;
wire [45:0] concat_7067;
wire [41:0] subW_3160;
wire [31:0] mul_3916;
wire [8:0] slice_4672;
wire [32:0] lsl_765;
wire [130:0] concat_5428;
wire [41:0] subW_1521;
wire [47:0] addW_6184;
wire [33:0] add_2277;
wire [34:0] addW_6940;
wire [13:0] slice_3033;
wire [7:0] slice_3789;
wire [16:0] mulnw_4545;
wire [34:0] addW_638;
wire [7:0] slice_5301;
wire [133:0] subW_1394;
wire [7:0] slice_6057;
wire [67:0] subW_2150;
wire [31:0] slice_6813;
wire [63:0] slice_2906;
wire [17:0] slice_7569;
wire [13:0] slice_3662;
wire [32:0] slice_4418;
wire [7:0] slice_511;
wire [19:0] addW_5174;
wire [15:0] slice_1267;
wire [35:0] mul_5930;
wire [31:0] slice_2023;
wire [66:0] concat_6686;
wire [19:0] addW_2779;
wire [19:0] addW_7442;
wire [15:0] mul_3535;
wire [31:0] slice_4291;
wire [34:0] addW_384;
wire [1029:0] concat_5047;
wire [31:0] slice_1140;
wire [25:0] lsl_5803;
wire [7:0] slice_1896;
wire [16:0] slice_6559;
wire [19:0] addW_2652;
wire [15:0] slice_7315;
wire [19:0] addW_3408;
wire [15:0] slice_4164;
wire [13:0] slice_257;
wire [71:0] subW_4920;
wire [7:0] slice_1013;
wire [31:0] mul_5676;
wire [17:0] slice_1769;
wire [64:0] slice_6432;
wire [51:0] addW_2525;
wire [66:0] addW_7188;
wire [7:0] slice_3281;
wire [15:0] slice_4037;
wire [13:0] slice_130;
wire [50:0] addW_4793;
wire [39:0] mul_886;
wire [17:0] add_5549;
wire [32:0] lsl_1642;
wire [32:0] lsl_6305;
wire [31:0] slice_2398;
wire [13:0] slice_7061;
wire [17:0] slice_3154;
wire [64:0] slice_3910;
wire [33:0] mul_4666;
wire [31:0] mul_759;
wire [15:0] slice_5422;
wire [17:0] slice_1515;
wire [45:0] concat_6178;
wire [7:0] slice_2271;
wire [15:0] mulnw_6934;
wire [33:0] add_3027;
wire [16:0] mulnw_3783;
wire [7:0] slice_4539;
wire [41:0] subW_632;
wire [7:0] slice_5295;
wire [70:0] subW_1388;
wire [7:0] slice_6051;
wire [26:0] add_2144;
wire [51:0] addW_6807;
wire [98:0] addW_2900;
wire [34:0] addW_7563;
wire [40:0] subW_3656;
wire [34:0] addW_4412;
wire [7:0] slice_505;
wire [17:0] slice_5168;
wire [33:0] addW_1261;
wire [13:0] slice_5924;
wire [39:0] mul_2017;
wire [15:0] mul_6680;
wire [17:0] slice_2773;
wire [27:0] mul_7436;
wire [7:0] slice_3529;
wire [31:0] slice_4285;
wire [15:0] mulnw_378;
wire [127:0] slice_5041;
wire [127:0] slice_1134;
wire [32:0] lsl_5797;
wire [16:0] mulnw_1890;
wire [47:0] addW_6553;
wire [17:0] slice_2646;
wire [32:0] slice_7309;
wire [17:0] slice_3402;
wire [50:0] addW_4158;
wire [33:0] add_251;
wire [40:0] subW_4914;
wire [8:0] slice_1007;
wire [31:0] slice_5670;
wire [34:0] addW_1763;
wire [195:0] addW_6426;
wire [49:0] concat_2519;
wire [68:0] subW_7182;
wire [16:0] mulnw_3275;
wire [97:0] concat_4031;
wire [130:0] concat_124;
wire [17:0] add_4787;
wire [17:0] slice_880;
wire [16:0] mulnw_5543;
wire [15:0] mul_1636;
wire [31:0] mul_6299;
wire [39:0] mul_2392;
wire [50:0] addW_7055;
wire [34:0] addW_3148;
wire [387:0] concat_3904;
wire [65:0] addW_4660;
wire [66:0] addW_753;
wire [25:0] lsl_5416;
wire [31:0] slice_1509;
wire [13:0] slice_6172;
wire [8:0] slice_2265;
wire [8:0] slice_6928;
wire [7:0] slice_3021;
wire [7:0] slice_3777;
wire [15:0] slice_4533;
wire [17:0] slice_626;
wire [16:0] mulnw_5289;
wire [39:0] mul_1382;
wire [16:0] mulnw_6045;
wire [16:0] mulnw_2138;
wire [49:0] concat_6801;
wire [34:0] addW_2894;
wire [15:0] slice_7557;
wire [35:0] mul_3650;
wire [15:0] mulnw_4406;
wire [16:0] mulnw_499;
wire [65:0] concat_5162;
wire [41:0] subW_1255;
wire [40:0] subW_5918;
wire [17:0] slice_2011;
wire [7:0] slice_6674;
wire [66:0] concat_2767;
wire [15:0] slice_7430;
wire [26:0] add_3523;
wire [51:0] addW_4279;
wire [8:0] slice_372;
wire [197:0] addW_5035;
wire [131:0] concat_1128;
wire [31:0] mul_5791;
wire [7:0] slice_1884;
wire [45:0] concat_6547;
wire [31:0] slice_2640;
wire [130:0] addW_7303;
wire [65:0] concat_3396;
wire [17:0] add_4152;
wire [7:0] slice_245;
wire [35:0] mul_4908;
wire [33:0] mul_1001;
wire [39:0] mul_5664;
wire [17:0] slice_1757;
wire [71:0] subW_6420;
wire [15:0] slice_2513;
wire [33:0] add_7176;
wire [7:0] slice_3269;
wire [40:0] subW_4025;
wire [15:0] slice_118;
wire [16:0] mulnw_4781;
wire [127:0] slice_874;
wire [25:0] lsl_5537;
wire [7:0] slice_1630;
wire [16:0] slice_6293;
wire [17:0] slice_2386;
wire [17:0] add_7049;
wire [17:0] slice_3142;
wire [132:0] subW_3898;
wire [68:0] subW_4654;
wire [195:0] concat_747;
wire [32:0] lsl_5410;
wire [41:0] subW_1503;
wire [63:0] slice_6166;
wire [33:0] mul_2259;
wire [17:0] add_6922;
wire [7:0] slice_3015;
wire [15:0] slice_3771;
wire [97:0] concat_4527;
wire [31:0] slice_620;
wire [7:0] slice_5283;
wire [17:0] slice_1376;
wire [7:0] slice_6039;
wire [33:0] add_2132;
wire [15:0] slice_6795;
wire [15:0] mulnw_2888;
wire [25:0] lsl_7551;
wire [63:0] slice_3644;
wire [8:0] slice_4400;
wire [7:0] slice_493;
wire [19:0] addW_5156;
wire [17:0] slice_1249;
wire [35:0] mul_5912;
wire [31:0] slice_2005;
wire [26:0] add_6668;
wire [15:0] mul_2761;
wire [25:0] lsl_7424;
wire [15:0] mulnw_3517;
wire [49:0] concat_4273;
wire [17:0] add_366;
wire [71:0] subW_5029;
wire [17:0] slice_1122;
wire [66:0] addW_5785;
wire [15:0] slice_1878;
wire [13:0] slice_6541;
wire [67:0] subW_2634;
wire [196:0] addW_7297;
wire [19:0] addW_3390;
wire [16:0] mulnw_4146;
wire [7:0] slice_239;
wire [15:0] slice_4902;
wire [31:0] slice_995;
wire [17:0] slice_5658;
wire [19:0] addW_1751;
wire [40:0] subW_6414;
wire [66:0] concat_2507;
wire [7:0] slice_7170;
wire [15:0] slice_3263;
wire [35:0] mul_4019;
wire [25:0] lsl_112;
wire [25:0] lsl_4775;
wire [255:0] slice_868;
wire [32:0] lsl_5531;
wire [15:0] slice_1624;
wire [47:0] addW_6287;
wire [31:0] slice_2380;
wire [16:0] mulnw_7043;
wire [19:0] addW_3136;
wire [69:0] concat_3892;
wire [33:0] add_4648;
wire [67:0] subW_741;
wire [15:0] mul_5404;
wire [17:0] slice_1497;
wire [132:0] subW_6160;
wire [32:0] slice_2253;
wire [16:0] mulnw_6916;
wire [16:0] mulnw_3009;
wire [97:0] concat_3765;
wire [40:0] subW_4521;
wire [34:0] addW_614;
wire [15:0] slice_5277;
wire [34:0] addW_1370;
wire [15:0] slice_6033;
wire [7:0] slice_2126;
wire [65:0] concat_6789;
wire [8:0] slice_2882;
wire [32:0] lsl_7545;
wire [259:0] concat_3638;
wire [17:0] add_4394;
wire [15:0] slice_487;
wire [17:0] slice_5150;
wire [31:0] slice_1243;
wire [63:0] slice_5906;
wire [39:0] mul_1999;
wire [15:0] mulnw_6662;
wire [7:0] slice_2755;
wire [32:0] lsl_7418;
wire [49:0] concat_3511;
wire [15:0] slice_4267;
wire [16:0] mulnw_360;
wire [40:0] subW_5023;
wire [19:0] addW_1116;
wire [131:0] concat_5779;
wire [32:0] slice_1872;
wire [47:0] addW_6535;
wire [26:0] add_2628;
wire [71:0] subW_7291;
wire [17:0] slice_3384;
wire [25:0] lsl_4140;
wire [16:0] mulnw_233;
wire [47:0] addW_4896;
wire [39:0] mul_989;
wire [31:0] slice_5652;
wire [27:0] mul_1745;
wire [35:0] mul_6408;
wire [15:0] mul_2501;
wire [7:0] slice_7164;
wire [32:0] slice_3257;
wire [13:0] slice_4013;
wire [32:0] lsl_106;
wire [32:0] lsl_4769;
wire [260:0] concat_862;
wire [31:0] mul_5525;
wire [32:0] slice_1618;
wire [45:0] concat_6281;
wire [26:0] add_2374;
wire [25:0] lsl_7037;
wire [27:0] mul_3130;
wire [19:0] addW_3886;
wire [7:0] slice_4642;
wire [26:0] add_735;
wire [7:0] slice_5398;
wire [31:0] slice_1491;
wire [69:0] concat_6154;
wire [127:0] slice_2247;
wire [15:0] slice_6910;
wire [7:0] slice_3003;
wire [40:0] subW_3759;
wire [35:0] mul_4515;
wire [15:0] mulnw_608;
wire [66:0] concat_5271;
wire [41:0] subW_1364;
wire [97:0] concat_6027;
wire [8:0] slice_2120;
wire [19:0] addW_6783;
wire [17:0] add_2876;
wire [15:0] mul_7539;
wire [31:0] slice_3632;
wire [16:0] mulnw_4388;
wire [32:0] slice_481;
wire [31:0] slice_5144;
wire [41:0] subW_1237;
wire [127:0] slice_5900;
wire [17:0] slice_1993;
wire [49:0] concat_6656;
wire [26:0] add_2749;
wire [15:0] mul_7412;
wire [16:0] slice_3505;
wire [65:0] concat_4261;
wire [15:0] slice_354;
wire [35:0] mul_5017;
wire [31:0] mul_1110;
wire [17:0] slice_5773;
wire [98:0] addW_1866;
wire [45:0] concat_6529;
wire [16:0] mulnw_2622;
wire [40:0] subW_7285;
wire [255:0] slice_3378;
wire [32:0] lsl_4134;
wire [7:0] slice_227;
wire [45:0] concat_4890;
wire [17:0] slice_983;
wire [26:0] add_5646;
wire [15:0] slice_1739;
wire [15:0] slice_6402;
wire [7:0] slice_2495;
wire [16:0] mulnw_7158;
wire [98:0] addW_3251;
wire [40:0] subW_4007;
wire [15:0] mul_100;
wire [31:0] mul_4763;
wire [32:0] slice_856;
wire [65:0] addW_5519;
wire [34:0] addW_1612;
wire [13:0] slice_6275;
wire [16:0] mulnw_2368;
wire [32:0] lsl_7031;
wire [15:0] slice_3124;
wire [17:0] slice_3880;
wire [7:0] slice_4636;
wire [16:0] mulnw_729;
wire [15:0] slice_5392;
wire [31:0] slice_1485;
wire [19:0] addW_6148;
wire [131:0] concat_2241;
wire [16:0] slice_6904;
wire [15:0] slice_2997;
wire [35:0] mul_3753;
wire [13:0] slice_4509;
wire [8:0] slice_602;
wire [15:0] mul_5265;
wire [17:0] slice_1358;
wire [40:0] subW_6021;
wire [33:0] mul_2114;
wire [17:0] slice_6777;
wire [16:0] mulnw_2870;
wire [7:0] slice_7533;
wire [51:0] addW_3626;
wire [15:0] slice_4382;
wire [98:0] addW_475;
wire [70:0] subW_5138;
wire [17:0] slice_1231;
wire [263:0] subW_5894;
wire [127:0] slice_1987;
wire [16:0] slice_6650;
wire [15:0] mulnw_2743;
wire [7:0] slice_7406;
wire [65:0] concat_3499;
wire [19:0] addW_4255;
wire [33:0] addW_348;
wire [15:0] slice_5011;
wire [31:0] slice_1104;
wire [19:0] addW_5767;
wire [34:0] addW_1860;
wire [13:0] slice_6523;
wire [33:0] add_2616;
wire [35:0] mul_7279;
wire [516:0] concat_3372;
wire [31:0] mul_4128;
wire [15:0] slice_221;
wire [13:0] slice_4884;
wire [31:0] slice_977;
wire [16:0] mulnw_5640;
wire [25:0] lsl_1733;
wire [47:0] addW_6396;
wire [26:0] add_2489;
wire [7:0] slice_7152;
wire [34:0] addW_3245;
wire [35:0] mul_4001;
wire [7:0] slice_94;
wire [64:0] slice_4757;
wire [51:0] addW_850;
wire [130:0] concat_5513;
wire [15:0] mulnw_1606;
wire [47:0] addW_6269;
wire [33:0] add_2362;
wire [31:0] mul_7025;
wire [25:0] lsl_3118;
wire [98:0] concat_3874;
wire [16:0] mulnw_4630;
wire [33:0] add_723;
wire [33:0] addW_5386;
wire [51:0] addW_1479;
wire [17:0] slice_6142;
wire [17:0] slice_2235;
wire [31:0] slice_6898;
wire [32:0] slice_2991;
wire [13:0] slice_3747;
wire [40:0] subW_4503;
wire [17:0] add_596;
wire [7:0] slice_5259;
wire [31:0] slice_1352;
wire [35:0] mul_6015;
wire [31:0] slice_2108;
wire [66:0] concat_6771;
wire [15:0] slice_2864;
wire [15:0] slice_7527;
wire [49:0] concat_3620;
wire [16:0] slice_4376;
wire [34:0] addW_469;
wire [39:0] mul_5132;
wire [31:0] slice_1225;
wire [133:0] concat_5888;
wire [63:0] slice_1981;
wire [50:0] addW_6644;
wire [49:0] concat_2737;
wire [15:0] slice_7400;
wire [19:0] addW_3493;
wire [17:0] slice_4249;
wire [41:0] subW_342;
wire [50:0] addW_5005;
wire [39:0] mul_1098;
wire [31:0] mul_5761;
wire [15:0] mulnw_1854;
wire [131:0] concat_6517;
wire [7:0] slice_2610;
wire [15:0] slice_7273;
wire [63:0] slice_3366;
wire [16:0] slice_4122;
wire [32:0] slice_215;
wire [50:0] addW_4878;
wire [39:0] mul_971;
wire [33:0] add_5634;
wire [32:0] lsl_1727;
wire [45:0] concat_6390;
wire [15:0] mulnw_2483;
wire [15:0] slice_7146;
wire [15:0] mulnw_3239;
wire [63:0] slice_3995;
wire [388:0] concat_4751;
wire [49:0] concat_844;
wire [15:0] slice_5507;
wire [8:0] slice_1600;
wire [45:0] concat_6263;
wire [7:0] slice_2356;
wire [64:0] slice_7019;
wire [32:0] lsl_3112;
wire [40:0] subW_3868;
wire [7:0] slice_4624;
wire [7:0] slice_717;
wire [17:0] slice_5380;
wire [49:0] concat_1473;
wire [98:0] concat_6136;
wire [19:0] addW_2229;
wire [50:0] addW_6892;
wire [98:0] addW_2985;
wire [40:0] subW_3741;
wire [35:0] mul_4497;
wire [16:0] mulnw_590;
wire [26:0] add_5253;
wire [34:0] addW_1346;
wire [13:0] slice_6009;
wire [39:0] mul_2102;
wire [15:0] mul_6765;
wire [33:0] addW_2858;
wire [32:0] slice_7521;
wire [15:0] slice_3614;
wire [31:0] slice_4370;
wire [15:0] mulnw_463;
wire [17:0] slice_5126;
wire [31:0] slice_1219;
wire [17:0] slice_5882;
wire [100:0] addW_1975;
wire [17:0] add_6638;
wire [16:0] slice_2731;
wire [32:0] slice_7394;
wire [17:0] slice_3487;
wire [66:0] concat_4243;
wire [17:0] slice_336;
wire [17:0] add_4999;
wire [17:0] slice_1092;
wire [31:0] slice_5755;
wire [8:0] slice_1848;
wire [17:0] slice_6511;
wire [8:0] slice_2604;
wire [50:0] addW_7267;
wire [100:0] addW_3360;
wire [33:0] add_4116;
wire [130:0] concat_209;
wire [17:0] add_4872;
wire [17:0] slice_965;
wire [7:0] slice_5628;
wire [15:0] mul_1721;
wire [13:0] slice_6384;
wire [49:0] concat_2477;
wire [97:0] concat_7140;
wire [8:0] slice_3233;
wire [99:0] addW_3989;
wire [15:0] slice_82;
wire [132:0] subW_4745;
wire [15:0] slice_838;
wire [25:0] lsl_5501;
wire [17:0] add_1594;
wire [13:0] slice_6257;
wire [8:0] slice_2350;
wire [260:0] concat_7013;
wire [15:0] mul_3106;
wire [35:0] mul_3862;
wire [15:0] slice_4618;
wire [8:0] slice_711;
wire [19:0] addW_5374;
wire [15:0] slice_1467;
wire [40:0] subW_6130;
wire [31:0] mul_2223;
wire [17:0] add_6886;
wire [34:0] addW_2979;
wire [35:0] mul_3735;
wire [63:0] slice_4491;
wire [15:0] slice_584;
wire [15:0] mulnw_5247;
wire [15:0] mulnw_1340;
wire [40:0] subW_6003;
wire [17:0] slice_2096;
wire [7:0] slice_6759;
wire [41:0] subW_2852;
wire [34:0] addW_7515;
wire [65:0] concat_3608;
wire [50:0] addW_4364;
wire [8:0] slice_457;
wire [34:0] addW_5120;
wire [50:0] addW_1213;
wire [19:0] addW_5876;
wire [41:0] subW_1969;
wire [16:0] mulnw_6632;
wire [194:0] concat_2725;
wire [31:0] slice_7388;
wire [65:0] concat_3481;
wire [15:0] mul_4237;
wire [31:0] slice_330;
wire [16:0] mulnw_4993;
wire [31:0] slice_1086;
wire [39:0] mul_5749;
wire [17:0] add_1842;
wire [19:0] addW_6505;
wire [33:0] mul_2598;
wire [17:0] add_7261;
wire [41:0] subW_3354;
wire [7:0] slice_4110;
wire [15:0] slice_203;
wire [16:0] mulnw_4866;
wire [13:0] slice_959;
wire [8:0] slice_5622;
wire [7:0] slice_1715;
wire [50:0] addW_6378;
wire [16:0] slice_2471;
wire [40:0] subW_7134;
wire [17:0] add_3227;
wire [41:0] subW_3983;
wire [69:0] concat_4739;
wire [32:0] slice_832;
wire [32:0] lsl_5495;
wire [16:0] mulnw_1588;
wire [130:0] concat_6251;
wire [33:0] mul_2344;
wire [32:0] slice_7007;
wire [7:0] slice_3100;
wire [13:0] slice_3856;
wire [97:0] concat_4612;
wire [33:0] mul_705;
wire [27:0] mul_5368;
wire [65:0] concat_1461;
wire [35:0] mul_6124;
wire [31:0] slice_2217;
wire [16:0] mulnw_6880;
wire [15:0] mulnw_2973;
wire [63:0] slice_3729;
wire [260:0] concat_4485;
wire [129:0] addW_578;
wire [49:0] concat_5241;
wire [8:0] slice_1334;
wire [35:0] mul_5997;
wire [31:0] slice_2090;
wire [26:0] add_6753;
wire [17:0] slice_2846;
wire [15:0] mulnw_7509;
wire [19:0] addW_3602;
wire [17:0] add_4358;
wire [17:0] add_451;
wire [41:0] subW_5114;
wire [17:0] add_1207;
wire [31:0] mul_5870;
wire [17:0] slice_1963;
wire [25:0] lsl_6626;
wire [67:0] subW_2719;
wire [51:0] addW_7382;
wire [19:0] addW_3475;
wire [7:0] slice_4231;
wire [41:0] subW_324;
wire [25:0] lsl_4987;
wire [26:0] add_1080;
wire [17:0] slice_5743;
wire [16:0] mulnw_1836;
wire [31:0] mul_6499;
wire [31:0] slice_2592;
wire [16:0] mulnw_7255;
wire [17:0] slice_3348;
wire [7:0] slice_4104;
wire [25:0] lsl_197;
wire [25:0] lsl_4860;
wire [68:0] subW_953;
wire [33:0] mul_5616;
wire [15:0] slice_1709;
wire [17:0] add_6372;
wire [50:0] addW_2465;
wire [35:0] mul_7128;
wire [16:0] mulnw_3221;
wire [17:0] slice_3977;
wire [31:0] slice_70;
wire [19:0] addW_4733;
wire [26:0] add_826;
wire [15:0] mul_5489;
wire [15:0] slice_1582;
wire [15:0] slice_6245;
wire [64:0] slice_2338;
wire [51:0] addW_7001;
wire [15:0] slice_3094;
wire [33:0] add_3850;
wire [40:0] subW_4606;
wire [31:0] slice_699;
wire [17:0] slice_5362;
wire [19:0] addW_1455;
wire [13:0] slice_6118;
wire [39:0] mul_2211;
wire [25:0] lsl_6874;
wire [8:0] slice_2967;
wire [98:0] addW_3723;
wire [32:0] slice_4479;
wire [16:0] slice_5235;
wire [17:0] add_1328;
wire [63:0] slice_5991;
wire [39:0] mul_2084;
wire [15:0] mulnw_6747;
wire [31:0] slice_2840;
wire [8:0] slice_7503;
wire [17:0] slice_3596;
wire [16:0] mulnw_4352;
wire [16:0] mulnw_445;
wire [17:0] slice_5108;
wire [16:0] mulnw_1201;
wire [32:0] slice_5864;
wire [34:0] addW_1957;
wire [32:0] lsl_6620;
wire [26:0] add_2713;
wire [49:0] concat_7376;
wire [17:0] slice_3469;
wire [26:0] add_4225;
wire [17:0] slice_318;
wire [32:0] lsl_4981;
wire [16:0] mulnw_1074;
wire [31:0] slice_5737;
wire [15:0] slice_1830;
wire [31:0] slice_6493;
wire [39:0] mul_2586;
wire [25:0] lsl_7249;
wire [34:0] addW_3342;
wire [16:0] mulnw_4098;
wire [32:0] lsl_191;
wire [32:0] lsl_4854;
wire [33:0] add_947;
wire [32:0] slice_5610;
wire [32:0] slice_1703;
wire [16:0] mulnw_6366;
wire [17:0] add_2459;
wire [13:0] slice_7122;
wire [15:0] slice_3215;
wire [34:0] addW_3971;
wire [39:0] mul_64;
wire [17:0] slice_4727;
wire [16:0] mulnw_820;
wire [7:0] slice_5483;
wire [16:0] slice_1576;
wire [25:0] lsl_6239;
wire [69:0] concat_2332;
wire [49:0] concat_6995;
wire [32:0] slice_3088;
wire [7:0] slice_3844;
wire [35:0] mul_4600;
wire [39:0] mul_693;
wire [19:0] addW_5356;
wire [17:0] slice_1449;
wire [33:0] add_6112;
wire [17:0] slice_2205;
wire [32:0] lsl_6868;
wire [17:0] add_2961;
wire [34:0] addW_3717;
wire [51:0] addW_4473;
wire [133:0] subW_566;
wire [195:0] concat_5229;
wire [16:0] mulnw_1322;
wire [98:0] addW_5985;
wire [17:0] slice_2078;
wire [49:0] concat_6741;
wire [41:0] subW_2834;
wire [17:0] add_7497;
wire [66:0] concat_3590;
wire [25:0] lsl_4346;
wire [15:0] slice_439;
wire [31:0] slice_5102;
wire [25:0] lsl_1195;
wire [26:0] add_5858;
wire [15:0] slice_1951;
wire [31:0] mul_6614;
wire [16:0] mulnw_2707;
wire [15:0] slice_7370;
wire [31:0] slice_3463;
wire [15:0] mulnw_4219;
wire [31:0] slice_312;
wire [31:0] mul_4975;
wire [33:0] add_1068;
wire [26:0] add_5731;
wire [33:0] addW_1824;
wire [39:0] mul_6487;
wire [17:0] slice_2580;
wire [32:0] lsl_7243;
wire [15:0] slice_3336;
wire [7:0] slice_4092;
wire [15:0] mul_185;
wire [31:0] mul_4848;
wire [7:0] slice_941;
wire [63:0] slice_5604;
wire [64:0] slice_1697;
wire [25:0] lsl_6360;
wire [16:0] mulnw_2453;
wire [40:0] subW_7116;
wire [33:0] addW_3209;
wire [17:0] slice_3965;
wire [17:0] slice_58;
wire [98:0] concat_4721;
wire [33:0] add_814;
wire [15:0] slice_5477;
wire [31:0] slice_1570;
wire [32:0] lsl_6233;
wire [19:0] addW_2326;
wire [15:0] slice_6989;
wire [129:0] addW_3082;
wire [7:0] slice_3838;
wire [13:0] slice_4594;
wire [17:0] slice_687;
wire [27:0] mul_5350;
wire [66:0] concat_1443;
wire [7:0] slice_6106;
wire [31:0] slice_2199;
wire [31:0] mul_6862;
wire [16:0] mulnw_2955;
wire [15:0] mulnw_3711;
wire [49:0] concat_4467;
wire [70:0] subW_560;
wire [67:0] subW_5223;
wire [15:0] slice_1316;
wire [34:0] addW_5979;
wire [13:0] slice_2072;
wire [16:0] slice_6735;
wire [17:0] slice_2828;
wire [16:0] mulnw_7491;
wire [15:0] mul_3584;
wire [32:0] lsl_4340;
wire [33:0] addW_433;
wire [34:0] addW_5096;
wire [32:0] lsl_1189;
wire [16:0] mulnw_5852;
wire [25:0] lsl_1945;
wire [66:0] addW_6608;
wire [33:0] add_2701;
wire [65:0] concat_7364;
wire [67:0] subW_3457;
wire [49:0] concat_4213;
wire [127:0] slice_306;
wire [16:0] slice_4969;
wire [7:0] slice_1062;
wire [16:0] mulnw_5725;
wire [41:0] subW_1818;
wire [17:0] slice_6481;
wire [31:0] slice_2574;
wire [31:0] mul_7237;
wire [25:0] lsl_3330;
wire [15:0] slice_4086;
wire [7:0] slice_179;
wire [64:0] slice_4842;
wire [7:0] slice_935;
wire [99:0] addW_5598;
wire [255:0] slice_1691;
wire [32:0] lsl_6354;
wire [25:0] lsl_2447;
wire [35:0] mul_7110;
wire [41:0] subW_3203;
wire [19:0] addW_3959;
wire [31:0] slice_52;
wire [40:0] subW_4715;
wire [7:0] slice_808;
wire [33:0] addW_5471;
wire [50:0] addW_1564;
wire [15:0] mul_6227;
wire [17:0] slice_2320;
wire [66:0] concat_6983;
wire [133:0] subW_3076;
wire [16:0] mulnw_3832;
wire [40:0] subW_4588;
wire [31:0] slice_681;
wire [31:0] slice_5344;
wire [15:0] mul_1437;
wire [7:0] slice_6100;
wire [26:0] add_2193;
wire [16:0] slice_6856;
wire [15:0] slice_2949;
wire [8:0] slice_3705;
wire [15:0] slice_4461;
wire [39:0] mul_554;
wire [26:0] add_5217;
wire [16:0] slice_1310;
wire [15:0] mulnw_5973;
wire [68:0] subW_2066;
wire [32:0] slice_6729;
wire [31:0] slice_2822;
wire [15:0] slice_7485;
wire [7:0] slice_3578;
wire [31:0] mul_4334;
wire [41:0] subW_427;
wire [15:0] mulnw_5090;
wire [31:0] mul_1183;
wire [33:0] add_5846;
wire [32:0] lsl_1939;
wire [130:0] concat_6602;
wire [7:0] slice_2695;
wire [19:0] addW_7358;
wire [26:0] add_3451;
wire [16:0] slice_4207;
wire [131:0] concat_300;
wire [33:0] add_4963;
wire [8:0] slice_1056;
wire [33:0] add_5719;
wire [17:0] slice_1812;
wire [31:0] slice_6475;
wire [39:0] mul_2568;
wire [16:0] slice_7231;
wire [32:0] lsl_3324;
wire [32:0] slice_4080;
wire [15:0] slice_173;
wire [99:0] addW_4836;
wire [16:0] mulnw_929;
wire [41:0] subW_5592;
wire [260:0] concat_1685;
wire [31:0] mul_6348;
wire [32:0] lsl_2441;
wire [63:0] slice_7104;
wire [17:0] slice_3197;
wire [27:0] mul_3953;
wire [39:0] mul_46;
wire [35:0] mul_4709;
wire [8:0] slice_802;
wire [17:0] slice_5465;
wire [17:0] add_1558;
wire [7:0] slice_6221;
wire [98:0] concat_2314;
wire [15:0] mul_6977;
wire [70:0] subW_3070;
wire [7:0] slice_3826;
wire [35:0] mul_4582;
wire [39:0] mul_675;
wire [135:0] subW_5338;
wire [7:0] slice_1431;
wire [16:0] mulnw_6094;
wire [16:0] mulnw_2187;
wire [47:0] addW_6850;
wire [33:0] addW_2943;
wire [17:0] add_3699;
wire [66:0] concat_4455;
wire [17:0] slice_548;
wire [16:0] mulnw_5211;
wire [31:0] slice_1304;
wire [8:0] slice_5967;
wire [33:0] add_2060;
wire [773:0] concat_6723;
wire [127:0] slice_2816;
wire [16:0] slice_7479;
wire [26:0] add_3572;
wire [16:0] slice_4328;
wire [17:0] slice_421;
wire [8:0] slice_5084;
wire [16:0] slice_1177;
wire [7:0] slice_5840;
wire [15:0] mul_1933;
wire [15:0] slice_6596;
wire [8:0] slice_2689;
wire [17:0] slice_7352;
wire [16:0] mulnw_3445;
wire [32:0] slice_4201;
wire [17:0] slice_294;
wire [7:0] slice_4957;
wire [33:0] mul_1050;
wire [7:0] slice_5713;
wire [31:0] slice_1806;
wire [26:0] add_6469;
wire [17:0] slice_2562;
wire [33:0] add_7225;
wire [15:0] mul_3318;
wire [98:0] addW_4074;
wire [33:0] addW_167;
wire [41:0] subW_4830;
wire [7:0] slice_923;
wire [17:0] slice_5586;
wire [32:0] slice_1679;
wire [65:0] addW_6342;
wire [31:0] mul_2435;
wire [99:0] addW_7098;
wire [31:0] slice_3191;
wire [15:0] slice_3947;
wire [17:0] slice_40;
wire [13:0] slice_4703;
wire [33:0] mul_796;
wire [19:0] addW_5459;
wire [16:0] mulnw_1552;
wire [15:0] slice_6215;
wire [40:0] subW_2308;
wire [7:0] slice_6971;
wire [39:0] mul_3064;
wire [15:0] slice_3820;
wire [63:0] slice_4576;
wire [17:0] slice_669;
wire [70:0] subW_5332;
wire [26:0] add_1425;
wire [7:0] slice_6088;
wire [33:0] add_2181;
wire [45:0] concat_6844;
wire [41:0] subW_2937;
wire [1032:0] subW_7600;
wire [16:0] mulnw_3693;
wire [15:0] mul_4449;
wire [34:0] addW_542;
wire [33:0] add_5205;
wire [50:0] addW_1298;
wire [17:0] add_5961;
wire [7:0] slice_2054;
wire [261:0] subW_6717;
wire [131:0] concat_2810;
wire [31:0] slice_7473;
wire [15:0] mulnw_3566;
wire [47:0] addW_4322;
wire [31:0] slice_415;
wire [17:0] add_5078;
wire [47:0] addW_1171;
wire [8:0] slice_5834;
wire [7:0] slice_1927;
wire [25:0] lsl_6590;
wire [33:0] mul_2683;
wire [66:0] concat_7346;
wire [33:0] add_3439;
wire [516:0] concat_4195;
wire [19:0] addW_288;
wire [7:0] slice_4951;
wire [65:0] addW_1044;
wire [8:0] slice_5707;
wire [41:0] subW_1800;
wire [16:0] mulnw_6463;
wire [127:0] slice_2556;
wire [7:0] slice_7219;
wire [7:0] slice_3312;
wire [34:0] addW_4068;
wire [17:0] slice_161;
wire [17:0] slice_4824;
wire [15:0] slice_917;
wire [34:0] addW_5580;
wire [51:0] addW_1673;
wire [130:0] concat_6336;
wire [66:0] addW_2429;
wire [41:0] subW_7092;
wire [41:0] subW_3185;
wire [25:0] lsl_3941;
wire [33:0] add_4697;
wire [15:0] slice_790;
wire [27:0] mul_5453;
wire [25:0] lsl_1546;
wire [33:0] addW_6209;
wire [35:0] mul_2302;
wire [26:0] add_6965;
wire [17:0] slice_3058;
wire [32:0] slice_3814;
wire [98:0] addW_4570;
wire [13:0] slice_663;
wire [39:0] mul_5326;
wire [15:0] mulnw_1419;
wire [15:0] slice_6082;
wire [7:0] slice_2175;
wire [13:0] slice_6838;
wire [17:0] slice_2931;
wire [520:0] subW_7594;
wire [15:0] slice_3687;
wire [7:0] slice_4443;
wire [41:0] subW_536;
wire [7:0] slice_5199;
wire [17:0] add_1292;
wire [16:0] mulnw_5955;
wire [7:0] slice_2048;
wire [133:0] concat_6711;
wire [17:0] slice_2804;
wire [51:0] addW_7467;
wire [49:0] concat_3560;
wire [45:0] concat_4316;
wire [41:0] subW_409;
wire [16:0] mulnw_5072;
wire [45:0] concat_1165;
wire [33:0] mul_5828;
wire [15:0] slice_1921;
wire [32:0] lsl_6584;
wire [31:0] slice_2677;
wire [15:0] mul_7340;
wire [7:0] slice_3433;
wire [63:0] slice_4189;
wire [31:0] mul_282;
wire [16:0] mulnw_4945;
wire [68:0] subW_1038;
wire [33:0] mul_5701;
wire [17:0] slice_1794;
wire [33:0] add_6457;
wire [127:0] slice_2550;
wire [7:0] slice_7213;
wire [15:0] slice_3306;
wire [15:0] mulnw_4062;
wire [19:0] addW_155;
wire [34:0] addW_4818;
wire [97:0] concat_911;
wire [17:0] slice_5574;
wire [49:0] concat_1667;
wire [15:0] slice_6330;
wire [64:0] slice_2423;
wire [17:0] slice_7086;
wire [17:0] slice_3179;
wire [32:0] lsl_3935;
wire [255:0] slice_28;
wire [7:0] slice_4691;
wire [25:0] lsl_784;
wire [17:0] slice_5447;
wire [32:0] lsl_1540;
wire [17:0] slice_6203;
wire [13:0] slice_2296;
wire [15:0] mulnw_6959;
wire [34:0] addW_3052;
wire [98:0] addW_3808;
wire [34:0] addW_4564;
wire [71:0] subW_657;
wire [17:0] slice_5320;
wire [49:0] concat_1413;
wire [32:0] slice_6076;
wire [8:0] slice_2169;
wire [47:0] addW_6832;
wire [31:0] slice_2925;
wire [262:0] concat_7588;
wire [33:0] addW_3681;
wire [26:0] add_4437;
wire [17:0] slice_530;
wire [8:0] slice_5193;
wire [16:0] mulnw_1286;
wire [15:0] slice_5949;
wire [16:0] mulnw_2042;
wire [17:0] slice_6705;
wire [19:0] addW_2798;
wire [49:0] concat_7461;
wire [16:0] slice_3554;
wire [13:0] slice_4310;
wire [17:0] slice_403;
wire [15:0] slice_5066;
wire [13:0] slice_1159;
wire [15:0] slice_5822;
wire [32:0] slice_1915;
wire [15:0] mul_6578;
wire [39:0] mul_2671;
wire [7:0] slice_7334;
wire [8:0] slice_3427;
wire [100:0] addW_4183;
wire [7:0] slice_4939;
wire [33:0] add_1032;
wire [64:0] slice_5695;
wire [31:0] slice_1788;
wire [7:0] slice_6451;
wire [519:0] subW_2544;
wire [16:0] mulnw_7207;
wire [32:0] slice_3300;
wire [8:0] slice_4056;
wire [27:0] mul_149;
wire [17:0] slice_4812;
wire [40:0] subW_905;
wire [19:0] addW_5568;
wire [15:0] slice_1661;
wire [25:0] lsl_6324;
wire [69:0] concat_2417;
wire [34:0] addW_7080;
wire [31:0] slice_3173;
wire [15:0] mul_3929;
wire [31:0] slice_22;
wire [7:0] slice_4685;
wire [32:0] lsl_778;
wire [19:0] addW_5441;
wire [31:0] mul_1534;
wire [19:0] addW_6197;
wire [33:0] add_2290;
wire [49:0] concat_6953;
wire [41:0] subW_3046;
wire [34:0] addW_3802;
wire [15:0] mulnw_4558;
wire [40:0] subW_651;
wire [34:0] addW_5314;
wire [16:0] slice_1407;
wire [98:0] addW_6070;
wire [33:0] mul_2163;
wire [45:0] concat_6826;
wire [41:0] subW_2919;
wire [32:0] slice_7582;
wire [41:0] subW_3675;
wire [15:0] mulnw_4431;
wire [31:0] slice_524;
wire [33:0] mul_5187;
wire [25:0] lsl_1280;
wire [33:0] addW_5943;
wire [7:0] slice_2036;
wire [19:0] addW_6699;
wire [31:0] mul_2792;
wire [15:0] slice_7455;
wire [194:0] concat_3548;
wire [47:0] addW_4304;
wire [31:0] slice_397;
wire [128:0] slice_5060;
wire [47:0] addW_1153;
wire [25:0] lsl_5816;
wire [34:0] addW_1909;
wire [7:0] slice_6572;
wire [17:0] slice_2665;
wire [26:0] add_7328;
wire [33:0] mul_3421;
wire [41:0] subW_4177;
wire [41:0] subW_270;
wire [15:0] slice_4933;
wire [7:0] slice_1026;
wire [69:0] concat_5689;
wire [31:0] slice_1782;
wire [8:0] slice_6445;
wire [263:0] subW_2538;
wire [7:0] slice_7201;
wire [34:0] addW_3294;
wire [17:0] add_4050;
wire [17:0] slice_143;
wire [19:0] addW_4806;
wire [35:0] mul_899;
wire [27:0] mul_5562;
wire [66:0] concat_1655;
wire [32:0] lsl_6318;
wire [19:0] addW_2411;
wire [17:0] slice_7074;
wire [31:0] slice_3167;
wire [7:0] slice_3923;
wire [127:0] slice_16;
wire [16:0] mulnw_4679;
wire [15:0] mul_772;
wire [27:0] mul_5435;
wire [16:0] slice_1528;
wire [27:0] mul_6191;
wire [7:0] slice_2284;
wire [16:0] slice_6947;
wire [17:0] slice_3040;
wire [15:0] mulnw_3796;
wire [8:0] slice_4552;
wire [35:0] mul_645;
wire [34:0] addW_5308;
wire [64:0] slice_1401;
wire [34:0] addW_6064;
wire [65:0] addW_2157;
wire [13:0] slice_6820;
wire [17:0] slice_2913;
wire [51:0] addW_7576;
wire [17:0] slice_3669;
wire [49:0] concat_4425;
wire [34:0] addW_518;
wire [31:0] slice_5181;
wire [32:0] lsl_1274;
wire [41:0] subW_5937;
wire [15:0] slice_2030;
wire [31:0] mul_6693;
wire [31:0] slice_2786;
wire [65:0] concat_7449;
wire [67:0] subW_3542;
wire [45:0] concat_4298;
wire [31:0] slice_391;
wire [128:0] slice_5054;
wire [45:0] concat_1147;
wire [32:0] lsl_5810;
wire [15:0] mulnw_1903;
wire [15:0] slice_6566;
wire [31:0] slice_2659;
wire [15:0] mulnw_7322;
wire [31:0] slice_3415;
wire [17:0] slice_4171;
wire [17:0] slice_264;
wire [32:0] slice_4927;
wire [7:0] slice_1020;
wire [19:0] addW_5683;
wire [51:0] addW_1776;
wire [33:0] mul_6439;
wire [133:0] concat_2532;
wire [15:0] slice_7195;
wire [15:0] mulnw_3288;
wire [16:0] mulnw_4044;
wire [19:0] addW_137;
wire [27:0] mul_4800;
wire [13:0] slice_893;
wire [15:0] slice_5556;
wire [15:0] mul_1649;
wire [15:0] mul_6312;
wire [17:0] slice_2405;
wire [19:0] addW_7068;
wire [51:0] addW_3161;
wire [15:0] slice_3917;
wire [511:0] slice_10;
wire [7:0] slice_4673;
wire [7:0] slice_766;
wire [63:0] slice_5429;
wire [47:0] addW_1522;
wire [17:0] slice_6185;
wire [7:0] slice_2278;
wire [50:0] addW_6941;
wire [31:0] slice_3034;
wire [8:0] slice_3790;
wire [17:0] add_4546;
wire [15:0] slice_639;
wire [15:0] mulnw_5302;
wire [195:0] addW_1395;
wire [15:0] mulnw_6058;
wire [68:0] subW_2151;
wire [131:0] concat_6814;
wire [31:0] slice_2907;
wire [49:0] concat_7570;
wire [31:0] slice_3663;
wire [16:0] slice_4419;
wire [15:0] mulnw_512;
wire [39:0] mul_5175;
wire [31:0] mul_1268;
wire [17:0] slice_5931;
wire [97:0] concat_2024;
wire [32:0] slice_6687;
wire [39:0] mul_2780;
wire [19:0] addW_7443;
wire [26:0] add_3536;
wire [13:0] slice_4292;
wire [50:0] addW_385;
wire [511:0] slice_5048;
wire [13:0] slice_1141;
wire [15:0] mul_5804;
wire [8:0] slice_1897;
wire [33:0] addW_6560;
wire [39:0] mul_2653;
wire [49:0] concat_7316;
wire [39:0] mul_3409;
wire [34:0] addW_4165;
wire [31:0] slice_258;
wire [99:0] addW_4921;
wire [16:0] mulnw_1014;
wire [17:0] slice_5677;
wire [49:0] concat_1770;
wire [32:0] slice_6433;
wire [17:0] slice_2526;
wire [32:0] slice_7189;
wire [8:0] slice_3282;
wire [15:0] slice_4038;
wire [27:0] mul_131;
wire [15:0] slice_4794;
wire [40:0] subW_887;
wire [25:0] lsl_5550;
wire [7:0] slice_1643;
wire [7:0] slice_6306;
wire [98:0] concat_2399;
wire [27:0] mul_7062;
wire [49:0] concat_3155;
wire [32:0] slice_3911;
wire [15:0] slice_4667;
wire [15:0] slice_760;
wire [66:0] concat_5423;
wire [45:0] concat_1516;
wire [19:0] addW_6179;
wire [16:0] mulnw_2272;
wire [17:0] add_6935;
wire [34:0] addW_3028;
wire [17:0] add_3784;
wire [16:0] mulnw_4540;
wire [47:0] addW_633;
wire [8:0] slice_5296;
wire [71:0] subW_1389;
wire [8:0] slice_6052;
wire [33:0] add_2145;
wire [17:0] slice_6808;
wire [31:0] slice_2901;
wire [15:0] slice_7564;
wire [41:0] subW_3657;
wire [50:0] addW_4413;
wire [8:0] slice_506;
wire [17:0] slice_5169;
wire [16:0] slice_1262;
wire [31:0] slice_5925;
wire [40:0] subW_2018;
wire [26:0] add_6681;
wire [17:0] slice_2774;
wire [17:0] slice_7437;
wire [16:0] mulnw_3530;
wire [131:0] concat_4286;
wire [17:0] add_379;
wire [517:0] concat_5042;
wire [63:0] slice_1135;
wire [7:0] slice_5798;
wire [17:0] add_1891;
wire [17:0] slice_6554;
wire [17:0] slice_2647;
wire [16:0] slice_7310;
wire [17:0] slice_3403;
wire [15:0] slice_4159;
wire [34:0] addW_252;
wire [41:0] subW_4915;
wire [7:0] slice_1008;
wire [98:0] concat_5671;
wire [15:0] slice_1764;
wire [63:0] slice_6427;
wire [19:0] addW_2520;
wire [98:0] addW_7183;
wire [17:0] add_3276;
wire [33:0] addW_4032;
wire [63:0] slice_125;
wire [25:0] lsl_4788;
wire [35:0] mul_881;
wire [32:0] lsl_5544;
wire [26:0] add_1637;
wire [15:0] slice_6300;
wire [40:0] subW_2393;
wire [15:0] slice_7056;
wire [15:0] slice_3149;
wire [129:0] addW_3905;
wire [32:0] slice_4661;
wire [32:0] slice_754;
wire [15:0] mul_5417;
wire [13:0] slice_1510;
wire [27:0] mul_6173;
wire [7:0] slice_2266;
wire [16:0] mulnw_6929;
wire [15:0] mulnw_3022;
wire [16:0] mulnw_3778;
wire [15:0] slice_4534;
wire [45:0] concat_627;
wire [17:0] add_5290;
wire [40:0] subW_1383;
wire [17:0] add_6046;
wire [7:0] slice_2139;
wire [19:0] addW_6802;
wire [50:0] addW_2895;
wire [66:0] concat_7558;
wire [17:0] slice_3651;
wire [17:0] add_4407;
wire [17:0] add_500;
wire [31:0] slice_5163;
wire [47:0] addW_1256;
wire [41:0] subW_5919;
wire [35:0] mul_2012;
wire [16:0] mulnw_6675;
wire [31:0] slice_2768;
wire [66:0] concat_7431;
wire [33:0] add_3524;
wire [17:0] slice_4280;
wire [16:0] mulnw_373;
wire [64:0] slice_5036;
wire [132:0] subW_1129;
wire [15:0] slice_5792;
wire [16:0] mulnw_1885;
wire [19:0] addW_6548;
wire [13:0] slice_2641;
wire [64:0] slice_7304;
wire [31:0] slice_3397;
wire [25:0] lsl_4153;
wire [15:0] mulnw_246;
wire [17:0] slice_4909;
wire [15:0] slice_1002;
wire [40:0] subW_5665;
wire [65:0] concat_1758;
wire [99:0] addW_6421;
wire [31:0] mul_2514;
wire [34:0] addW_7177;
wire [16:0] mulnw_3270;
wire [41:0] subW_4026;
wire [66:0] concat_119;
wire [32:0] lsl_4782;
wire [63:0] slice_875;
wire [15:0] mul_5538;
wire [15:0] mulnw_1631;
wire [33:0] addW_6294;
wire [35:0] mul_2387;
wire [25:0] lsl_7050;
wire [65:0] concat_3143;
wire [133:0] subW_3899;
wire [98:0] addW_4655;
wire [7:0] slice_5411;
wire [47:0] addW_1504;
wire [31:0] slice_6167;
wire [15:0] slice_2260;
wire [25:0] lsl_6923;
wire [8:0] slice_3016;
wire [15:0] slice_3772;
wire [33:0] addW_4528;
wire [13:0] slice_621;
wire [16:0] mulnw_5284;
wire [35:0] mul_1377;
wire [16:0] mulnw_6040;
wire [7:0] slice_2133;
wire [31:0] mul_6796;
wire [17:0] add_2889;
wire [15:0] mul_7552;
wire [31:0] slice_3645;
wire [16:0] mulnw_4401;
wire [16:0] mulnw_494;
wire [39:0] mul_5157;
wire [45:0] concat_1250;
wire [17:0] slice_5913;
wire [13:0] slice_2006;
wire [33:0] add_6669;
wire [26:0] add_2762;
wire [15:0] mul_7425;
wire [7:0] slice_3518;
wire [19:0] addW_4274;
wire [25:0] lsl_367;
wire [100:0] addW_5030;
wire [69:0] concat_1123;
wire [32:0] slice_5786;
wire [15:0] slice_1879;
wire [27:0] mul_6542;
wire [68:0] subW_2635;
wire [63:0] slice_7298;
wire [39:0] mul_3391;
wire [32:0] lsl_4147;
wire [8:0] slice_240;
wire [34:0] addW_4903;
wire [97:0] concat_996;
wire [35:0] mul_5659;
wire [19:0] addW_1752;
wire [41:0] subW_6415;
wire [32:0] slice_2508;
wire [15:0] mulnw_7171;
wire [15:0] slice_3264;
wire [17:0] slice_4020;
wire [15:0] mul_113;
wire [15:0] mul_4776;
wire [127:0] slice_869;
wire [7:0] slice_5532;
wire [49:0] concat_1625;
wire [17:0] slice_6288;
wire [13:0] slice_2381;
wire [32:0] lsl_7044;
wire [19:0] addW_3137;
wire [70:0] subW_3893;
wire [34:0] addW_4649;
wire [68:0] subW_742;
wire [26:0] add_5405;
wire [45:0] concat_1498;
wire [133:0] subW_6161;
wire [16:0] slice_2254;
wire [32:0] lsl_6917;
wire [17:0] add_3010;
wire [33:0] addW_3766;
wire [41:0] subW_4522;
wire [50:0] addW_615;
wire [15:0] slice_5278;
wire [15:0] slice_1371;
wire [15:0] slice_6034;
wire [16:0] mulnw_2127;
wire [31:0] slice_6790;
wire [16:0] mulnw_2883;
wire [7:0] slice_7546;
wire [127:0] slice_3639;
wire [25:0] lsl_4395;
wire [15:0] slice_488;
wire [17:0] slice_5151;
wire [13:0] slice_1244;
wire [31:0] slice_5907;
wire [40:0] subW_2000;
wire [7:0] slice_6663;
wire [16:0] mulnw_2756;
wire [7:0] slice_7419;
wire [8:0] slice_3512;
wire [31:0] mul_4268;
wire [32:0] lsl_361;
wire [41:0] subW_5024;
wire [19:0] addW_1117;
wire [64:0] slice_5780;
wire [16:0] slice_1873;
wire [17:0] slice_6536;
wire [33:0] add_2629;
wire [100:0] addW_7292;
wire [17:0] slice_3385;
wire [15:0] mul_4141;
wire [17:0] add_234;
wire [17:0] slice_4897;
wire [40:0] subW_990;
wire [13:0] slice_5653;
wire [17:0] slice_1746;
wire [17:0] slice_6409;
wire [26:0] add_2502;
wire [8:0] slice_7165;
wire [16:0] slice_3258;
wire [31:0] slice_4014;
wire [7:0] slice_107;
wire [7:0] slice_4770;
wire [261:0] subW_863;
wire [15:0] slice_5526;
wire [16:0] slice_1619;
wire [19:0] addW_6282;
wire [33:0] add_2375;
wire [15:0] mul_7038;
wire [17:0] slice_3131;
wire [39:0] mul_3887;
wire [15:0] mulnw_4643;
wire [33:0] add_736;
wire [15:0] mulnw_5399;
wire [13:0] slice_1492;
wire [70:0] subW_6155;
wire [388:0] concat_2248;
wire [31:0] mul_6911;
wire [16:0] mulnw_3004;
wire [41:0] subW_3760;
wire [17:0] slice_4516;
wire [17:0] add_609;
wire [32:0] slice_5272;
wire [47:0] addW_1365;
wire [33:0] addW_6028;
wire [7:0] slice_2121;
wire [39:0] mul_6784;
wire [25:0] lsl_2877;
wire [26:0] add_7540;
wire [131:0] concat_3633;
wire [32:0] lsl_4389;
wire [16:0] slice_482;
wire [13:0] slice_5145;
wire [47:0] addW_1238;
wire [63:0] slice_5901;
wire [35:0] mul_1994;
wire [8:0] slice_6657;
wire [33:0] add_2750;
wire [26:0] add_7413;
wire [33:0] mul_3506;
wire [31:0] slice_4262;
wire [31:0] mul_355;
wire [17:0] slice_5018;
wire [17:0] slice_1111;
wire [69:0] concat_5774;
wire [31:0] slice_1867;
wire [19:0] addW_6530;
wire [7:0] slice_2623;
wire [41:0] subW_7286;
wire [127:0] slice_3379;
wire [7:0] slice_4135;
wire [16:0] mulnw_228;
wire [19:0] addW_4891;
wire [35:0] mul_984;
wire [33:0] add_5647;
wire [66:0] concat_1740;
wire [34:0] addW_6403;
wire [16:0] mulnw_2496;
wire [17:0] add_7159;
wire [31:0] slice_3252;
wire [41:0] subW_4008;
wire [26:0] add_101;
wire [15:0] slice_4764;
wire [133:0] concat_857;
wire [32:0] slice_5520;
wire [50:0] addW_1613;
wire [27:0] mul_6276;
wire [7:0] slice_2369;
wire [7:0] slice_7032;
wire [66:0] concat_3125;
wire [17:0] slice_3881;
wire [8:0] slice_4637;
wire [7:0] slice_730;
wire [49:0] concat_5393;
wire [131:0] concat_1486;
wire [39:0] mul_6149;
wire [132:0] subW_2242;
wire [66:0] addW_6905;
wire [15:0] slice_2998;
wire [17:0] slice_3754;
wire [31:0] slice_4510;
wire [16:0] mulnw_603;
wire [26:0] add_5266;
wire [45:0] concat_1359;
wire [41:0] subW_6022;
wire [15:0] slice_2115;
wire [17:0] slice_6778;
wire [32:0] lsl_2871;
wire [15:0] mulnw_7534;
wire [17:0] slice_3627;
wire [31:0] mul_4383;
wire [31:0] slice_476;
wire [71:0] subW_5139;
wire [45:0] concat_1232;
wire [264:0] subW_5895;
wire [63:0] slice_1988;
wire [33:0] mul_6651;
wire [7:0] slice_2744;
wire [15:0] mulnw_7407;
wire [31:0] slice_3500;
wire [39:0] mul_4256;
wire [16:0] slice_349;
wire [34:0] addW_5012;
wire [98:0] concat_1105;
wire [19:0] addW_5768;
wire [50:0] addW_1861;
wire [27:0] mul_6524;
wire [7:0] slice_2617;
wire [17:0] slice_7280;
wire [255:0] slice_3373;
wire [15:0] slice_4129;
wire [15:0] slice_222;
wire [27:0] mul_4885;
wire [13:0] slice_978;
wire [7:0] slice_5641;
wire [15:0] mul_1734;
wire [17:0] slice_6397;
wire [33:0] add_2490;
wire [16:0] mulnw_7153;
wire [50:0] addW_3246;
wire [17:0] slice_4002;
wire [15:0] mulnw_95;
wire [32:0] slice_4758;
wire [17:0] slice_851;
wire [63:0] slice_5514;
wire [17:0] add_1607;
wire [17:0] slice_6270;
wire [7:0] slice_2363;
wire [15:0] slice_7026;
wire [15:0] mul_3119;
wire [34:0] addW_3875;
wire [17:0] add_4631;
wire [7:0] slice_724;
wire [16:0] slice_5387;
wire [17:0] slice_1480;
wire [17:0] slice_6143;
wire [69:0] concat_2236;
wire [130:0] concat_6899;
wire [16:0] slice_2992;
wire [31:0] slice_3748;
wire [41:0] subW_4504;
wire [25:0] lsl_597;
wire [16:0] mulnw_5260;
wire [13:0] slice_1353;
wire [17:0] slice_6016;
wire [97:0] concat_2109;
wire [31:0] slice_6772;
wire [31:0] mul_2865;
wire [49:0] concat_7528;
wire [19:0] addW_3621;
wire [66:0] addW_4377;
wire [50:0] addW_470;
wire [40:0] subW_5133;
wire [13:0] slice_1226;
wire [134:0] subW_5889;
wire [260:0] concat_1982;
wire [15:0] slice_6645;
wire [8:0] slice_2738;
wire [49:0] concat_7401;
wire [39:0] mul_3494;
wire [17:0] slice_4250;
wire [47:0] addW_343;
wire [15:0] slice_5006;
wire [40:0] subW_1099;
wire [17:0] slice_5762;
wire [17:0] add_1855;
wire [63:0] slice_6518;
wire [16:0] mulnw_2611;
wire [34:0] addW_7274;
wire [260:0] concat_3367;
wire [32:0] slice_4123;
wire [16:0] slice_216;
wire [15:0] slice_4879;
wire [40:0] subW_972;
wire [7:0] slice_5635;
wire [7:0] slice_1728;
wire [19:0] addW_6391;
wire [7:0] slice_2484;
wire [15:0] slice_7147;
wire [17:0] add_3240;
wire [31:0] slice_3996;
wire [8:0] slice_89;
wire [130:0] addW_4752;
wire [19:0] addW_845;
wire [66:0] concat_5508;
wire [16:0] mulnw_1601;
wire [19:0] addW_6264;
wire [16:0] mulnw_2357;
wire [32:0] slice_7020;
wire [7:0] slice_3113;
wire [41:0] subW_3869;
wire [16:0] mulnw_4625;
wire [16:0] mulnw_718;
wire [65:0] concat_5381;
wire [19:0] addW_1474;
wire [34:0] addW_6137;
wire [19:0] addW_2230;
wire [15:0] slice_6893;
wire [31:0] slice_2986;
wire [41:0] subW_3742;
wire [17:0] slice_4498;
wire [32:0] lsl_591;
wire [33:0] add_5254;
wire [50:0] addW_1347;
wire [31:0] slice_6010;
wire [40:0] subW_2103;
wire [26:0] add_6766;
wire [16:0] slice_2859;
wire [16:0] slice_7522;
wire [31:0] mul_3615;
wire [130:0] concat_4371;
wire [17:0] add_464;
wire [35:0] mul_5127;
wire [130:0] concat_1220;
wire [69:0] concat_5883;
wire [32:0] slice_1976;
wire [25:0] lsl_6639;
wire [33:0] mul_2732;
wire [16:0] slice_7395;
wire [17:0] slice_3488;
wire [31:0] slice_4244;
wire [45:0] concat_337;
wire [25:0] lsl_5000;
wire [35:0] mul_1093;
wire [98:0] concat_5756;
wire [16:0] mulnw_1849;
wire [69:0] concat_6512;
wire [7:0] slice_2605;
wire [15:0] slice_7268;
wire [32:0] slice_3361;
wire [34:0] addW_4117;
wire [63:0] slice_210;
wire [25:0] lsl_4873;
wire [35:0] mul_966;
wire [16:0] mulnw_5629;
wire [26:0] add_1722;
wire [27:0] mul_6385;
wire [8:0] slice_2478;
wire [33:0] addW_7141;
wire [16:0] mulnw_3234;
wire [31:0] slice_3990;
wire [15:0] slice_83;
wire [133:0] subW_4746;
wire [31:0] mul_839;
wire [15:0] mul_5502;
wire [25:0] lsl_1595;
wire [27:0] mul_6258;
wire [7:0] slice_2351;
wire [128:0] slice_7014;
wire [26:0] add_3107;
wire [17:0] slice_3863;
wire [15:0] slice_4619;
wire [7:0] slice_712;
wire [19:0] addW_5375;
wire [31:0] mul_1468;
wire [41:0] subW_6131;
wire [17:0] slice_2224;
wire [25:0] lsl_6887;
wire [50:0] addW_2980;
wire [17:0] slice_3736;
wire [31:0] slice_4492;
wire [31:0] mul_585;
wire [7:0] slice_5248;
wire [17:0] add_1341;
wire [41:0] subW_6004;
wire [35:0] mul_2097;
wire [16:0] mulnw_6760;
wire [47:0] addW_2853;
wire [50:0] addW_7516;
wire [31:0] slice_3609;
wire [15:0] slice_4365;
wire [16:0] mulnw_458;
wire [15:0] slice_5121;
wire [15:0] slice_1214;
wire [19:0] addW_5877;
wire [51:0] addW_1970;
wire [32:0] lsl_6633;
wire [65:0] addW_2726;
wire [131:0] concat_7389;
wire [31:0] slice_3482;
wire [26:0] add_4238;
wire [13:0] slice_331;
wire [32:0] lsl_4994;
wire [13:0] slice_1087;
wire [40:0] subW_5750;
wire [25:0] lsl_1843;
wire [19:0] addW_6506;
wire [15:0] slice_2599;
wire [25:0] lsl_7262;
wire [51:0] addW_3355;
wire [15:0] mulnw_4111;
wire [66:0] concat_204;
wire [32:0] lsl_4867;
wire [63:0] slice_960;
wire [7:0] slice_5623;
wire [15:0] mulnw_1716;
wire [15:0] slice_6379;
wire [33:0] mul_2472;
wire [41:0] subW_7135;
wire [25:0] lsl_3228;
wire [51:0] addW_3984;
wire [16:0] slice_77;
wire [70:0] subW_4740;
wire [99:0] concat_833;
wire [7:0] slice_5496;
wire [32:0] lsl_1589;
wire [63:0] slice_6252;
wire [15:0] slice_2345;
wire [133:0] concat_7008;
wire [15:0] mulnw_3101;
wire [31:0] slice_3857;
wire [33:0] addW_4613;
wire [15:0] slice_706;
wire [17:0] slice_5369;
wire [31:0] slice_1462;
wire [17:0] slice_6125;
wire [98:0] concat_2218;
wire [32:0] lsl_6881;
wire [17:0] add_2974;
wire [31:0] slice_3730;
wire [127:0] slice_4486;
wire [64:0] slice_579;
wire [8:0] slice_5242;
wire [16:0] mulnw_1335;
wire [17:0] slice_5998;
wire [13:0] slice_2091;
wire [33:0] add_6754;
wire [45:0] concat_2847;
wire [17:0] add_7510;
wire [39:0] mul_3603;
wire [25:0] lsl_4359;
wire [25:0] lsl_452;
wire [47:0] addW_5115;
wire [25:0] lsl_1208;
wire [17:0] slice_5871;
wire [49:0] concat_1964;
wire [15:0] mul_6627;
wire [68:0] subW_2720;
wire [17:0] slice_7383;
wire [39:0] mul_3476;
wire [16:0] mulnw_4232;
wire [47:0] addW_325;
wire [15:0] mul_4988;
wire [33:0] add_1081;
wire [35:0] mul_5744;
wire [32:0] lsl_1837;
wire [17:0] slice_6500;
wire [97:0] concat_2593;
wire [32:0] lsl_7256;
wire [49:0] concat_3349;
wire [8:0] slice_4105;
wire [15:0] mul_198;
wire [15:0] mul_4861;
wire [98:0] addW_954;
wire [15:0] slice_5617;
wire [49:0] concat_1710;
wire [25:0] lsl_6373;
wire [15:0] slice_2466;
wire [17:0] slice_7129;
wire [32:0] lsl_3222;
wire [49:0] concat_3978;
wire [97:0] concat_71;
wire [39:0] mul_4734;
wire [33:0] add_827;
wire [26:0] add_5490;
wire [31:0] mul_1583;
wire [66:0] concat_6246;
wire [32:0] slice_2339;
wire [17:0] slice_7002;
wire [49:0] concat_3095;
wire [34:0] addW_3851;
wire [41:0] subW_4607;
wire [97:0] concat_700;
wire [65:0] concat_5363;
wire [39:0] mul_1456;
wire [31:0] slice_6119;
wire [40:0] subW_2212;
wire [15:0] mul_6875;
wire [16:0] mulnw_2968;
wire [31:0] slice_3724;
wire [133:0] concat_4480;
wire [33:0] mul_5236;
wire [25:0] lsl_1329;
wire [31:0] slice_5992;
wire [40:0] subW_2085;
wire [7:0] slice_6748;
wire [13:0] slice_2841;
wire [16:0] mulnw_7504;
wire [17:0] slice_3597;
wire [32:0] lsl_4353;
wire [32:0] lsl_446;
wire [45:0] concat_5109;
wire [32:0] lsl_1202;
wire [99:0] concat_5865;
wire [15:0] slice_1958;
wire [7:0] slice_6621;
wire [33:0] add_2714;
wire [19:0] addW_7377;
wire [17:0] slice_3470;
wire [33:0] add_4226;
wire [45:0] concat_319;
wire [7:0] slice_4982;
wire [7:0] slice_1075;
wire [13:0] slice_5738;
wire [31:0] mul_1831;
wire [98:0] concat_6494;
wire [40:0] subW_2587;
wire [15:0] mul_7250;
wire [15:0] slice_3343;
wire [17:0] add_4099;
wire [7:0] slice_192;
wire [7:0] slice_4855;
wire [34:0] addW_948;
wire [16:0] slice_5611;
wire [16:0] slice_1704;
wire [32:0] lsl_6367;
wire [25:0] lsl_2460;
wire [31:0] slice_7123;
wire [31:0] mul_3216;
wire [15:0] slice_3972;
wire [40:0] subW_65;
wire [17:0] slice_4728;
wire [7:0] slice_821;
wire [15:0] mulnw_5484;
wire [66:0] addW_1577;
wire [15:0] mul_6240;
wire [70:0] subW_2333;
wire [19:0] addW_6996;
wire [16:0] slice_3089;
wire [15:0] mulnw_3845;
wire [17:0] slice_4601;
wire [40:0] subW_694;
wire [19:0] addW_5357;
wire [17:0] slice_1450;
wire [34:0] addW_6113;
wire [35:0] mul_2206;
wire [7:0] slice_6869;
wire [25:0] lsl_2962;
wire [50:0] addW_3718;
wire [17:0] slice_4474;
wire [195:0] addW_567;
wire [66:0] addW_5230;
wire [32:0] lsl_1323;
wire [31:0] slice_5986;
wire [35:0] mul_2079;
wire [8:0] slice_6742;
wire [47:0] addW_2835;
wire [25:0] lsl_7498;
wire [31:0] slice_3591;
wire [15:0] mul_4347;
wire [31:0] mul_440;
wire [13:0] slice_5103;
wire [15:0] mul_1196;
wire [33:0] add_5859;
wire [66:0] concat_1952;
wire [15:0] slice_6615;
wire [7:0] slice_2708;
wire [31:0] mul_7371;
wire [13:0] slice_3464;
wire [7:0] slice_4220;
wire [13:0] slice_313;
wire [15:0] slice_4976;
wire [7:0] slice_1069;
wire [33:0] add_5732;
wire [16:0] slice_1825;
wire [40:0] subW_6488;
wire [35:0] mul_2581;
wire [7:0] slice_7244;
wire [66:0] concat_3337;
wire [16:0] mulnw_4093;
wire [26:0] add_186;
wire [15:0] slice_4849;
wire [15:0] mulnw_942;
wire [259:0] concat_5605;
wire [32:0] slice_1698;
wire [15:0] mul_6361;
wire [32:0] lsl_2454;
wire [41:0] subW_7117;
wire [16:0] slice_3210;
wire [65:0] concat_3966;
wire [35:0] mul_59;
wire [34:0] addW_4722;
wire [7:0] slice_815;
wire [49:0] concat_5478;
wire [130:0] concat_1571;
wire [7:0] slice_6234;
wire [39:0] mul_2327;
wire [31:0] mul_6990;
wire [64:0] slice_3083;
wire [8:0] slice_3839;
wire [31:0] slice_4595;
wire [35:0] mul_688;
wire [17:0] slice_5351;
wire [31:0] slice_1444;
wire [15:0] mulnw_6107;
wire [13:0] slice_2200;
wire [15:0] slice_6863;
wire [32:0] lsl_2956;
wire [17:0] add_3712;
wire [19:0] addW_4468;
wire [71:0] subW_561;
wire [68:0] subW_5224;
wire [31:0] mul_1317;
wire [50:0] addW_5980;
wire [63:0] slice_2073;
wire [33:0] mul_6736;
wire [45:0] concat_2829;
wire [32:0] lsl_7492;
wire [26:0] add_3585;
wire [7:0] slice_4341;
wire [16:0] slice_434;
wire [50:0] addW_5097;
wire [7:0] slice_1190;
wire [7:0] slice_5853;
wire [15:0] mul_1946;
wire [32:0] slice_6609;
wire [7:0] slice_2702;
wire [31:0] slice_7365;
wire [68:0] subW_3458;
wire [8:0] slice_4214;
wire [63:0] slice_307;
wire [32:0] slice_4970;
wire [16:0] mulnw_1063;
wire [7:0] slice_5726;
wire [47:0] addW_1819;
wire [35:0] mul_6482;
wire [13:0] slice_2575;
wire [15:0] slice_7238;
wire [15:0] mul_3331;
wire [15:0] slice_4087;
wire [15:0] mulnw_180;
wire [32:0] slice_4843;
wire [8:0] slice_936;
wire [31:0] slice_5599;
wire [772:0] concat_1692;
wire [7:0] slice_6355;
wire [15:0] mul_2448;
wire [17:0] slice_7111;
wire [47:0] addW_3204;
wire [19:0] addW_3960;
wire [13:0] slice_53;
wire [41:0] subW_4716;
wire [16:0] mulnw_809;
wire [16:0] slice_5472;
wire [15:0] slice_1565;
wire [26:0] add_6228;
wire [17:0] slice_2321;
wire [32:0] slice_6984;
wire [195:0] addW_3077;
wire [17:0] add_3833;
wire [41:0] subW_4589;
wire [13:0] slice_682;
wire [13:0] slice_5345;
wire [26:0] add_1438;
wire [8:0] slice_6101;
wire [33:0] add_2194;
wire [33:0] addW_6857;
wire [31:0] mul_2950;
wire [16:0] mulnw_3706;
wire [31:0] mul_4462;
wire [40:0] subW_555;
wire [33:0] add_5218;
wire [65:0] addW_1311;
wire [17:0] add_5974;
wire [98:0] addW_2067;
wire [16:0] slice_6730;
wire [13:0] slice_2823;
wire [31:0] mul_7486;
wire [16:0] mulnw_3579;
wire [15:0] slice_4335;
wire [47:0] addW_428;
wire [17:0] add_5091;
wire [15:0] slice_1184;
wire [7:0] slice_5847;
wire [7:0] slice_1940;
wire [63:0] slice_6603;
wire [16:0] mulnw_2696;
wire [39:0] mul_7359;
wire [33:0] add_3452;
wire [33:0] mul_4208;
wire [132:0] subW_301;
wire [34:0] addW_4964;
wire [7:0] slice_1057;
wire [7:0] slice_5720;
wire [45:0] concat_1813;
wire [13:0] slice_6476;
wire [40:0] subW_2569;
wire [32:0] slice_7232;
wire [7:0] slice_3325;
wire [16:0] slice_4081;
wire [49:0] concat_174;
wire [31:0] slice_4837;
wire [17:0] add_930;
wire [51:0] addW_5593;
wire [261:0] subW_1686;
wire [15:0] slice_6349;
wire [7:0] slice_2442;
wire [31:0] slice_7105;
wire [45:0] concat_3198;
wire [17:0] slice_3954;
wire [40:0] subW_47;
wire [17:0] slice_4710;
wire [7:0] slice_803;
wire [65:0] concat_5466;
wire [25:0] lsl_1559;
wire [15:0] mulnw_6222;
wire [34:0] addW_2315;
wire [26:0] add_6978;
wire [71:0] subW_3071;
wire [16:0] mulnw_3827;
wire [17:0] slice_4583;
wire [40:0] subW_676;
wire [196:0] addW_5339;
wire [16:0] mulnw_1432;
wire [17:0] add_6095;
wire [7:0] slice_2188;
wire [17:0] slice_6851;
wire [16:0] slice_2944;
wire [25:0] lsl_3700;
wire [32:0] slice_4456;
wire [35:0] mul_549;
wire [7:0] slice_5212;
wire [130:0] concat_1305;
wire [16:0] mulnw_5968;
wire [34:0] addW_2061;
wire [63:0] slice_2817;
wire [66:0] addW_7480;
wire [33:0] add_3573;
wire [33:0] addW_4329;
wire [45:0] concat_422;
wire [16:0] mulnw_5085;
wire [33:0] addW_1178;
wire [16:0] mulnw_5841;
wire [26:0] add_1934;
wire [66:0] concat_6597;
wire [7:0] slice_2690;
wire [17:0] slice_7353;
wire [7:0] slice_3446;
wire [16:0] slice_4202;
wire [69:0] concat_295;
wire [15:0] mulnw_4958;
wire [15:0] slice_1051;
wire [16:0] mulnw_5714;
wire [13:0] slice_1807;
wire [33:0] add_6470;
wire [35:0] mul_2563;
wire [34:0] addW_7226;
wire [26:0] add_3319;
wire [31:0] slice_4075;
wire [16:0] slice_168;
wire [51:0] addW_4831;
wire [16:0] mulnw_924;
wire [49:0] concat_5587;
wire [133:0] concat_1680;
wire [32:0] slice_6343;
wire [15:0] slice_2436;
wire [31:0] slice_7099;
wire [13:0] slice_3192;
wire [66:0] concat_3948;
wire [45:0] concat_41;
wire [31:0] slice_4704;
wire [15:0] slice_797;
wire [19:0] addW_5460;
wire [32:0] lsl_1553;
wire [49:0] concat_6216;
wire [41:0] subW_2309;
wire [16:0] mulnw_6972;
wire [40:0] subW_3065;
wire [15:0] slice_3821;
wire [31:0] slice_4577;
wire [35:0] mul_670;
wire [71:0] subW_5333;
wire [33:0] add_1426;
wire [16:0] mulnw_6089;
wire [7:0] slice_2182;
wire [19:0] addW_6845;
wire [47:0] addW_2938;
wire [1542:0] addW_7601;
wire [32:0] lsl_3694;
wire [26:0] add_4450;
wire [15:0] slice_543;
wire [7:0] slice_5206;
wire [15:0] slice_1299;
wire [25:0] lsl_5962;
wire [15:0] mulnw_2055;
wire [262:0] subW_6718;
wire [132:0] subW_2811;
wire [131:0] concat_7474;
wire [7:0] slice_3567;
wire [17:0] slice_4323;
wire [13:0] slice_416;
wire [25:0] lsl_5079;
wire [17:0] slice_1172;
wire [7:0] slice_5835;
wire [15:0] mulnw_1928;
wire [15:0] mul_6591;
wire [15:0] slice_2684;
wire [31:0] slice_7347;
wire [7:0] slice_3440;
wire [255:0] slice_4196;
wire [19:0] addW_289;
wire [8:0] slice_4952;
wire [32:0] slice_1045;
wire [7:0] slice_5708;
wire [47:0] addW_1801;
wire [7:0] slice_6464;
wire [63:0] slice_2557;
wire [15:0] mulnw_7220;
wire [15:0] mulnw_3313;
wire [50:0] addW_4069;
wire [65:0] concat_162;
wire [49:0] concat_4825;
wire [15:0] slice_918;
wire [15:0] slice_5581;
wire [17:0] slice_1674;
wire [63:0] slice_6337;
wire [32:0] slice_2430;
wire [51:0] addW_7093;
wire [47:0] addW_3186;
wire [15:0] mul_3942;
wire [34:0] addW_4698;
wire [66:0] concat_791;
wire [17:0] slice_5454;
wire [15:0] mul_1547;
wire [16:0] slice_6210;
wire [17:0] slice_2303;
wire [33:0] add_6966;
wire [35:0] mul_3059;
wire [16:0] slice_3815;
wire [31:0] slice_4571;
wire [63:0] slice_664;
wire [40:0] subW_5327;
wire [7:0] slice_1420;
wire [15:0] slice_6083;
wire [16:0] mulnw_2176;
wire [27:0] mul_6839;
wire [45:0] concat_2932;
wire [521:0] subW_7595;
wire [31:0] mul_3688;
wire [16:0] mulnw_4444;
wire [47:0] addW_537;
wire [16:0] mulnw_5200;
wire [25:0] lsl_1293;
wire [32:0] lsl_5956;
wire [8:0] slice_2049;
wire [134:0] subW_6712;
wire [69:0] concat_2805;
wire [17:0] slice_7468;
wire [8:0] slice_3561;
wire [19:0] addW_4317;
wire [47:0] addW_410;
wire [32:0] lsl_5073;
wire [19:0] addW_1166;
wire [15:0] slice_5829;
wire [49:0] concat_1922;
wire [7:0] slice_6585;
wire [97:0] concat_2678;
wire [26:0] add_7341;
wire [16:0] mulnw_3434;
wire [260:0] concat_4190;
wire [17:0] slice_283;
wire [17:0] add_4946;
wire [98:0] addW_1039;
wire [15:0] slice_5702;
wire [45:0] concat_1795;
wire [7:0] slice_6458;
wire [63:0] slice_2551;
wire [8:0] slice_7214;
wire [49:0] concat_3307;
wire [17:0] add_4063;
wire [19:0] addW_156;
wire [15:0] slice_4819;
wire [33:0] addW_912;
wire [65:0] concat_5575;
wire [19:0] addW_1668;
wire [66:0] concat_6331;
wire [196:0] concat_2424;
wire [49:0] concat_7087;
wire [45:0] concat_3180;
wire [7:0] slice_3936;
wire [127:0] slice_29;
wire [15:0] mulnw_4692;
wire [15:0] mul_785;
wire [65:0] concat_5448;
wire [7:0] slice_1541;
wire [65:0] concat_6204;
wire [31:0] slice_2297;
wire [7:0] slice_6960;
wire [15:0] slice_3053;
wire [31:0] slice_3809;
wire [50:0] addW_4565;
wire [99:0] addW_658;
wire [35:0] mul_5321;
wire [8:0] slice_1414;
wire [16:0] slice_6077;
wire [7:0] slice_2170;
wire [17:0] slice_6833;
wire [13:0] slice_2926;
wire [263:0] subW_7589;
wire [16:0] slice_3682;
wire [33:0] add_4438;
wire [45:0] concat_531;
wire [7:0] slice_5194;
wire [32:0] lsl_1287;
wire [31:0] mul_5950;
wire [17:0] add_2043;
wire [69:0] concat_6706;
wire [19:0] addW_2799;
wire [19:0] addW_7462;
wire [33:0] mul_3555;
wire [27:0] mul_4311;
wire [45:0] concat_404;
wire [31:0] mul_5067;
wire [27:0] mul_1160;
wire [66:0] concat_5823;
wire [16:0] slice_1916;
wire [26:0] add_6579;
wire [40:0] subW_2672;
wire [16:0] mulnw_7335;
wire [7:0] slice_3428;
wire [32:0] slice_4184;
wire [16:0] mulnw_4940;
wire [34:0] addW_1033;
wire [32:0] slice_5696;
wire [13:0] slice_1789;
wire [16:0] mulnw_6452;
wire [773:0] addW_2545;
wire [17:0] add_7208;
wire [16:0] slice_3301;
wire [16:0] mulnw_4057;
wire [17:0] slice_150;
wire [65:0] concat_4813;
wire [41:0] subW_906;
wire [19:0] addW_5569;
wire [31:0] mul_1662;
wire [15:0] mul_6325;
wire [70:0] subW_2418;
wire [15:0] slice_7081;
wire [13:0] slice_3174;
wire [26:0] add_3930;
wire [8:0] slice_4686;
wire [7:0] slice_779;
wire [19:0] addW_5442;
wire [15:0] slice_1535;
wire [19:0] addW_6198;
wire [34:0] addW_2291;
wire [8:0] slice_6954;
wire [47:0] addW_3047;
wire [50:0] addW_3803;
wire [17:0] add_4559;
wire [41:0] subW_652;
wire [15:0] slice_5315;
wire [33:0] mul_1408;
wire [31:0] slice_6071;
wire [15:0] slice_2164;
wire [19:0] addW_6827;
wire [47:0] addW_2920;
wire [133:0] concat_7583;
wire [47:0] addW_3676;
wire [7:0] slice_4432;
wire [13:0] slice_525;
wire [15:0] slice_5188;
wire [15:0] mul_1281;
wire [16:0] slice_5944;
wire [16:0] mulnw_2037;
wire [19:0] addW_6700;
wire [17:0] slice_2793;
wire [31:0] mul_7456;
wire [65:0] addW_3549;
wire [17:0] slice_4305;
wire [13:0] slice_398;
wire [64:0] slice_5061;
wire [17:0] slice_1154;
wire [15:0] mul_5817;
wire [50:0] addW_1910;
wire [15:0] mulnw_6573;
wire [35:0] mul_2666;
wire [33:0] add_7329;
wire [15:0] slice_3422;
wire [51:0] addW_4178;
wire [47:0] addW_271;
wire [15:0] slice_4934;
wire [15:0] mulnw_1027;
wire [70:0] subW_5690;
wire [131:0] concat_1783;
wire [7:0] slice_6446;
wire [264:0] subW_2539;
wire [16:0] mulnw_7202;
wire [50:0] addW_3295;
wire [25:0] lsl_4051;
wire [65:0] concat_144;
wire [19:0] addW_4807;
wire [17:0] slice_900;
wire [17:0] slice_5563;
wire [32:0] slice_1656;
wire [7:0] slice_6319;
wire [39:0] mul_2412;
wire [65:0] concat_7075;
wire [131:0] concat_3168;
wire [15:0] mulnw_3924;
wire [17:0] add_4680;
wire [26:0] add_773;
wire [17:0] slice_5436;
wire [33:0] addW_1529;
wire [17:0] slice_6192;
wire [15:0] mulnw_2285;
wire [33:0] mul_6948;
wire [45:0] concat_3041;
wire [17:0] add_3797;
wire [16:0] mulnw_4553;
wire [17:0] slice_646;
wire [50:0] addW_5309;
wire [32:0] slice_1402;
wire [50:0] addW_6065;
wire [32:0] slice_2158;
wire [27:0] mul_6821;
wire [45:0] concat_2914;
wire [17:0] slice_7577;
wire [45:0] concat_3670;
wire [8:0] slice_4426;
wire [50:0] addW_519;
wire [97:0] concat_5182;
wire [7:0] slice_1275;
wire [47:0] addW_5938;
wire [15:0] slice_2031;
wire [17:0] slice_6694;
wire [98:0] concat_2787;
wire [31:0] slice_7450;
wire [68:0] subW_3543;
wire [19:0] addW_4299;
wire [130:0] concat_392;
wire [64:0] slice_5055;
wire [19:0] addW_1148;
wire [7:0] slice_5811;
wire [17:0] add_1904;
wire [49:0] concat_6567;
wire [13:0] slice_2660;
wire [7:0] slice_7323;
wire [97:0] concat_3416;
wire [49:0] concat_4172;
wire [45:0] concat_265;
wire [16:0] slice_4928;
wire [8:0] slice_1021;
wire [39:0] mul_5684;
wire [17:0] slice_1777;
wire [15:0] slice_6440;
wire [134:0] subW_2533;
wire [15:0] slice_7196;
wire [17:0] add_3289;
wire [32:0] lsl_4045;
wire [19:0] addW_138;
wire [17:0] slice_4801;
wire [31:0] slice_894;
wire [66:0] concat_5557;
wire [26:0] add_1650;
wire [26:0] add_6313;
wire [17:0] slice_2406;
wire [19:0] addW_7069;
wire [17:0] slice_3162;
wire [49:0] concat_3918;
wire [16:0] mulnw_4674;
wire [15:0] mulnw_767;
wire [31:0] slice_5430;
wire [17:0] slice_1523;
wire [65:0] concat_6186;
wire [8:0] slice_2279;
wire [15:0] slice_6942;
wire [13:0] slice_3035;
wire [16:0] mulnw_3791;
wire [25:0] lsl_4547;
wire [34:0] addW_640;
wire [17:0] add_5303;
wire [63:0] slice_1396;
wire [17:0] add_6059;
wire [98:0] addW_2152;
wire [63:0] slice_6815;
wire [13:0] slice_2908;
wire [19:0] addW_7571;
wire [13:0] slice_3664;
wire [33:0] mul_4420;
wire [17:0] add_513;
wire [40:0] subW_5176;
wire [15:0] slice_1269;
wire [45:0] concat_5932;
wire [33:0] addW_2025;
wire [99:0] concat_6688;
wire [40:0] subW_2781;
wire [39:0] mul_7444;
wire [33:0] add_3537;
wire [27:0] mul_4293;
wire [15:0] slice_386;
wire [1541:0] concat_5049;
wire [27:0] mul_1142;
wire [26:0] add_5805;
wire [16:0] mulnw_1898;
wire [16:0] slice_6561;
wire [40:0] subW_2654;
wire [8:0] slice_7317;
wire [40:0] subW_3410;
wire [15:0] slice_4166;
wire [13:0] slice_259;
wire [31:0] slice_4922;
wire [17:0] add_1015;
wire [17:0] slice_5678;
wire [19:0] addW_1771;
wire [16:0] slice_6434;
wire [69:0] concat_2527;
wire [16:0] slice_7190;
wire [16:0] mulnw_3283;
wire [31:0] mul_4039;
wire [17:0] slice_132;
wire [66:0] concat_4795;
wire [41:0] subW_888;
wire [15:0] mul_5551;
wire [16:0] mulnw_1644;
wire [15:0] mulnw_6307;
wire [34:0] addW_2400;
wire [17:0] slice_7063;
wire [19:0] addW_3156;
wire [16:0] slice_3912;
wire [15:0] slice_4668;
wire [49:0] concat_761;
wire [67:0] subW_5424;
wire [19:0] addW_1517;
wire [19:0] addW_6180;
wire [17:0] add_2273;
wire [25:0] lsl_6936;
wire [50:0] addW_3029;
wire [25:0] lsl_3785;
wire [32:0] lsl_4541;
wire [17:0] slice_634;
wire [16:0] mulnw_5297;
wire [99:0] addW_1390;
wire [16:0] mulnw_6053;
wire [34:0] addW_2146;
wire [69:0] concat_6809;
wire [130:0] concat_2902;
wire [31:0] mul_7565;
wire [47:0] addW_3658;
wire [15:0] slice_4414;
wire [16:0] mulnw_507;
wire [35:0] mul_5170;
wire [33:0] addW_1263;
wire [13:0] slice_5926;
wire [41:0] subW_2019;
wire [33:0] add_6682;
wire [35:0] mul_2775;
wire [17:0] slice_7438;
wire [7:0] slice_3531;
wire [63:0] slice_4287;
wire [25:0] lsl_380;
wire [518:0] subW_5043;
wire [31:0] slice_1136;
wire [15:0] mulnw_5799;
wire [25:0] lsl_1892;
wire [65:0] concat_6555;
wire [35:0] mul_2648;
wire [33:0] mul_7311;
wire [35:0] mul_3404;
wire [66:0] concat_4160;
wire [50:0] addW_253;
wire [51:0] addW_4916;
wire [16:0] mulnw_1009;
wire [34:0] addW_5672;
wire [31:0] mul_1765;
wire [259:0] concat_6428;
wire [19:0] addW_2521;
wire [31:0] slice_7184;
wire [25:0] lsl_3277;
wire [16:0] slice_4033;
wire [31:0] slice_126;
wire [15:0] mul_4789;
wire [17:0] slice_882;
wire [7:0] slice_5545;
wire [33:0] add_1638;
wire [49:0] concat_6301;
wire [41:0] subW_2394;
wire [66:0] concat_7057;
wire [31:0] mul_3150;
wire [64:0] slice_3906;
wire [16:0] slice_4662;
wire [16:0] slice_755;
wire [26:0] add_5418;
wire [27:0] mul_1511;
wire [17:0] slice_6174;
wire [16:0] mulnw_2267;
wire [32:0] lsl_6930;
wire [17:0] add_3023;
wire [32:0] lsl_3779;
wire [31:0] mul_4535;
wire [19:0] addW_628;
wire [25:0] lsl_5291;
wire [41:0] subW_1384;
wire [25:0] lsl_6047;
wire [15:0] mulnw_2140;
wire [19:0] addW_6803;
wire [15:0] slice_2896;
wire [32:0] slice_7559;
wire [45:0] concat_3652;
wire [25:0] lsl_4408;
wire [25:0] lsl_501;
wire [13:0] slice_5164;
wire [17:0] slice_1257;
wire [47:0] addW_5920;
wire [17:0] slice_2013;
wire [7:0] slice_6676;
wire [13:0] slice_2769;
wire [31:0] slice_7432;
wire [7:0] slice_3525;
wire [69:0] concat_4281;
wire [32:0] lsl_374;
wire [262:0] concat_5037;
wire [133:0] subW_1130;
wire [49:0] concat_5793;
wire [32:0] lsl_1886;
wire [19:0] addW_6549;
wire [63:0] slice_2642;
wire [32:0] slice_7305;
wire [13:0] slice_3398;
wire [15:0] mul_4154;
wire [17:0] add_247;
wire [49:0] concat_4910;
wire [15:0] slice_1003;
wire [41:0] subW_5666;
wire [31:0] slice_1759;
wire [31:0] slice_6422;
wire [17:0] slice_2515;
wire [50:0] addW_7178;
wire [32:0] lsl_3271;
wire [47:0] addW_4027;
wire [67:0] subW_120;
wire [7:0] slice_4783;
wire [31:0] slice_876;
wire [26:0] add_5539;
wire [7:0] slice_1632;
wire [16:0] slice_6295;
wire [17:0] slice_2388;
wire [15:0] mul_7051;
wire [31:0] slice_3144;
wire [195:0] addW_3900;
wire [31:0] slice_4656;
wire [16:0] mulnw_5412;
wire [17:0] slice_1505;
wire [13:0] slice_6168;
wire [15:0] slice_2261;
wire [15:0] mul_6924;
wire [16:0] mulnw_3017;
wire [31:0] mul_3773;
wire [16:0] slice_4529;
wire [27:0] mul_622;
wire [32:0] lsl_5285;
wire [17:0] slice_1378;
wire [32:0] lsl_6041;
wire [8:0] slice_2134;
wire [17:0] slice_6797;
wire [25:0] lsl_2890;
wire [26:0] add_7553;
wire [13:0] slice_3646;
wire [32:0] lsl_4402;
wire [32:0] lsl_495;
wire [40:0] subW_5158;
wire [19:0] addW_1251;
wire [45:0] concat_5914;
wire [31:0] slice_2007;
wire [7:0] slice_6670;
wire [33:0] add_2763;
wire [26:0] add_7426;
wire [16:0] mulnw_3519;
wire [19:0] addW_4275;
wire [15:0] mul_368;
wire [32:0] slice_5031;
wire [70:0] subW_1124;
wire [16:0] slice_5787;
wire [31:0] mul_1880;
wire [17:0] slice_6543;
wire [98:0] addW_2636;
wire [260:0] concat_7299;
wire [40:0] subW_3392;
wire [7:0] slice_4148;
wire [16:0] mulnw_241;
wire [15:0] slice_4904;
wire [33:0] addW_997;
wire [17:0] slice_5660;
wire [39:0] mul_1753;
wire [51:0] addW_6416;
wire [99:0] concat_2509;
wire [17:0] add_7172;
wire [31:0] mul_3265;
wire [45:0] concat_4021;
wire [26:0] add_114;
wire [26:0] add_4777;
wire [63:0] slice_870;
wire [15:0] mulnw_5533;
wire [8:0] slice_1626;
wire [65:0] concat_6289;
wire [31:0] slice_2382;
wire [7:0] slice_7045;
wire [39:0] mul_3138;
wire [71:0] subW_3894;
wire [50:0] addW_4650;
wire [98:0] addW_743;
wire [33:0] add_5406;
wire [19:0] addW_1499;
wire [195:0] addW_6162;
wire [130:0] addW_2255;
wire [7:0] slice_6918;
wire [25:0] lsl_3011;
wire [16:0] slice_3767;
wire [47:0] addW_4523;
wire [15:0] slice_616;
wire [31:0] mul_5279;
wire [34:0] addW_1372;
wire [31:0] mul_6035;
wire [17:0] add_2128;
wire [98:0] concat_6791;
wire [32:0] lsl_2884;
wire [16:0] mulnw_7547;
wire [63:0] slice_3640;
wire [15:0] mul_4396;
wire [31:0] mul_489;
wire [35:0] mul_5152;
wire [27:0] mul_1245;
wire [13:0] slice_5908;
wire [41:0] subW_2001;
wire [16:0] mulnw_6664;
wire [7:0] slice_2757;
wire [16:0] mulnw_7420;
wire [7:0] slice_3513;
wire [17:0] slice_4269;
wire [7:0] slice_362;
wire [51:0] addW_5025;
wire [39:0] mul_1118;
wire [196:0] concat_5781;
wire [66:0] addW_1874;
wire [65:0] concat_6537;
wire [34:0] addW_2630;
wire [32:0] slice_7293;
wire [35:0] mul_3386;
wire [26:0] add_4142;
wire [25:0] lsl_235;
wire [65:0] concat_4898;
wire [41:0] subW_991;
wire [31:0] slice_5654;
wire [17:0] slice_1747;
wire [49:0] concat_6410;
wire [33:0] add_2503;
wire [16:0] mulnw_7166;
wire [66:0] addW_3259;
wire [13:0] slice_4015;
wire [16:0] mulnw_108;
wire [15:0] mulnw_4771;
wire [262:0] subW_864;
wire [49:0] concat_5527;
wire [33:0] mul_1620;
wire [19:0] addW_6283;
wire [34:0] addW_2376;
wire [26:0] add_7039;
wire [17:0] slice_3132;
wire [40:0] subW_3888;
wire [17:0] add_4644;
wire [34:0] addW_737;
wire [7:0] slice_5400;
wire [27:0] mul_1493;
wire [71:0] subW_6156;
wire [15:0] slice_6912;
wire [32:0] lsl_3005;
wire [47:0] addW_3761;
wire [45:0] concat_4517;
wire [25:0] lsl_610;
wire [16:0] slice_5273;
wire [17:0] slice_1366;
wire [16:0] slice_6029;
wire [16:0] mulnw_2122;
wire [40:0] subW_6785;
wire [15:0] mul_2878;
wire [33:0] add_7541;
wire [132:0] subW_3634;
wire [7:0] slice_4390;
wire [65:0] addW_483;
wire [63:0] slice_5146;
wire [17:0] slice_1239;
wire [31:0] slice_5902;
wire [17:0] slice_1995;
wire [7:0] slice_6658;
wire [7:0] slice_2751;
wire [33:0] add_7414;
wire [15:0] slice_3507;
wire [98:0] concat_4263;
wire [15:0] slice_356;
wire [49:0] concat_5019;
wire [17:0] slice_1112;
wire [70:0] subW_5775;
wire [130:0] concat_1868;
wire [19:0] addW_6531;
wire [15:0] mulnw_2624;
wire [51:0] addW_7287;
wire [63:0] slice_3380;
wire [15:0] mulnw_4136;
wire [32:0] lsl_229;
wire [19:0] addW_4892;
wire [17:0] slice_985;
wire [34:0] addW_5648;
wire [31:0] slice_1741;
wire [15:0] slice_6404;
wire [7:0] slice_2497;
wire [25:0] lsl_7160;
wire [130:0] concat_3253;
wire [47:0] addW_4009;
wire [33:0] add_102;
wire [49:0] concat_4765;
wire [134:0] subW_858;
wire [16:0] slice_5521;
wire [15:0] slice_1614;
wire [17:0] slice_6277;
wire [15:0] mulnw_2370;
wire [15:0] mulnw_7033;
wire [31:0] slice_3126;
wire [35:0] mul_3882;
wire [16:0] mulnw_4638;
wire [15:0] mulnw_731;
wire [8:0] slice_5394;
wire [63:0] slice_1487;
wire [40:0] subW_6150;
wire [133:0] subW_2243;
wire [32:0] slice_6906;
wire [31:0] mul_2999;
wire [45:0] concat_3755;
wire [13:0] slice_4511;
wire [32:0] lsl_604;
wire [33:0] add_5267;
wire [19:0] addW_1360;
wire [47:0] addW_6023;
wire [15:0] slice_2116;
wire [35:0] mul_6779;
wire [7:0] slice_2872;
wire [7:0] slice_7535;
wire [69:0] concat_3628;
wire [15:0] slice_4384;
wire [130:0] concat_477;
wire [99:0] addW_5140;
wire [19:0] addW_1233;
wire [389:0] addW_5896;
wire [31:0] slice_1989;
wire [15:0] slice_6652;
wire [16:0] mulnw_2745;
wire [7:0] slice_7408;
wire [97:0] concat_3501;
wire [40:0] subW_4257;
wire [33:0] addW_350;
wire [15:0] slice_5013;
wire [34:0] addW_1106;
wire [39:0] mul_5769;
wire [15:0] slice_1862;
wire [17:0] slice_6525;
wire [8:0] slice_2618;
wire [49:0] concat_7281;
wire [127:0] slice_3374;
wire [49:0] concat_4130;
wire [31:0] mul_223;
wire [17:0] slice_4886;
wire [31:0] slice_979;
wire [15:0] mulnw_5642;
wire [26:0] add_1735;
wire [65:0] concat_6398;
wire [7:0] slice_2491;
wire [32:0] lsl_7154;
wire [15:0] slice_3247;
wire [45:0] concat_4003;
wire [7:0] slice_96;
wire [16:0] slice_4759;
wire [69:0] concat_852;
wire [194:0] concat_5515;
wire [25:0] lsl_1608;
wire [65:0] concat_6271;
wire [8:0] slice_2364;
wire [49:0] concat_7027;
wire [26:0] add_3120;
wire [15:0] slice_3876;
wire [25:0] lsl_4632;
wire [8:0] slice_725;
wire [33:0] mul_5388;
wire [69:0] concat_1481;
wire [35:0] mul_6144;
wire [70:0] subW_2237;
wire [63:0] slice_6900;
wire [65:0] addW_2993;
wire [13:0] slice_3749;
wire [47:0] addW_4505;
wire [15:0] mul_598;
wire [7:0] slice_5261;
wire [27:0] mul_1354;
wire [45:0] concat_6017;
wire [33:0] addW_2110;
wire [13:0] slice_6773;
wire [15:0] slice_2866;
wire [8:0] slice_7529;
wire [19:0] addW_3622;
wire [32:0] slice_4378;
wire [15:0] slice_471;
wire [41:0] subW_5134;
wire [27:0] mul_1227;
wire [135:0] subW_5890;
wire [127:0] slice_1983;
wire [66:0] concat_6646;
wire [7:0] slice_2739;
wire [8:0] slice_7402;
wire [40:0] subW_3495;
wire [35:0] mul_4251;
wire [17:0] slice_344;
wire [66:0] concat_5007;
wire [41:0] subW_1100;
wire [17:0] slice_5763;
wire [25:0] lsl_1856;
wire [31:0] slice_6519;
wire [17:0] add_2612;
wire [15:0] slice_7275;
wire [261:0] subW_3368;
wire [16:0] slice_4124;
wire [65:0] addW_217;
wire [66:0] concat_4880;
wire [41:0] subW_973;
wire [8:0] slice_5636;
wire [16:0] mulnw_1729;
wire [19:0] addW_6392;
wire [16:0] mulnw_2485;
wire [31:0] mul_7148;
wire [25:0] lsl_3241;
wire [13:0] slice_3997;
wire [7:0] slice_90;
wire [64:0] slice_4753;
wire [19:0] addW_846;
wire [67:0] subW_5509;
wire [32:0] lsl_1602;
wire [19:0] addW_6265;
wire [17:0] add_2358;
wire [16:0] slice_7021;
wire [16:0] mulnw_3114;
wire [47:0] addW_3870;
wire [32:0] lsl_4626;
wire [17:0] add_719;
wire [31:0] slice_5382;
wire [19:0] addW_1475;
wire [15:0] slice_6138;
wire [39:0] mul_2231;
wire [66:0] concat_6894;
wire [130:0] concat_2987;
wire [47:0] addW_3743;
wire [45:0] concat_4499;
wire [7:0] slice_592;
wire [7:0] slice_5255;
wire [15:0] slice_1348;
wire [13:0] slice_6011;
wire [41:0] subW_2104;
wire [33:0] add_6767;
wire [33:0] addW_2860;
wire [33:0] mul_7523;
wire [17:0] slice_3616;
wire [63:0] slice_4372;
wire [25:0] lsl_465;
wire [17:0] slice_5128;
wire [63:0] slice_1221;
wire [70:0] subW_5884;
wire [133:0] concat_1977;
wire [15:0] mul_6640;
wire [15:0] slice_2733;
wire [33:0] mul_7396;
wire [35:0] mul_3489;
wire [13:0] slice_4245;
wire [19:0] addW_338;
wire [15:0] mul_5001;
wire [17:0] slice_1094;
wire [34:0] addW_5757;
wire [32:0] lsl_1850;
wire [70:0] subW_6513;
wire [16:0] mulnw_2606;
wire [66:0] concat_7269;
wire [133:0] concat_3362;
wire [50:0] addW_4118;
wire [194:0] concat_211;
wire [15:0] mul_4874;
wire [17:0] slice_967;
wire [17:0] add_5630;
wire [33:0] add_1723;
wire [17:0] slice_6386;
wire [7:0] slice_2479;
wire [16:0] slice_7142;
wire [32:0] lsl_3235;
wire [131:0] concat_3991;
wire [31:0] mul_84;
wire [195:0] addW_4747;
wire [17:0] slice_840;
wire [26:0] add_5503;
wire [15:0] mul_1596;
wire [17:0] slice_6259;
wire [16:0] mulnw_2352;
wire [64:0] slice_7015;
wire [33:0] add_3108;
wire [45:0] concat_3864;
wire [31:0] mul_4620;
wire [16:0] mulnw_713;
wire [39:0] mul_5376;
wire [17:0] slice_1469;
wire [47:0] addW_6132;
wire [17:0] slice_2225;
wire [15:0] mul_6888;
wire [15:0] slice_2981;
wire [45:0] concat_3737;
wire [13:0] slice_4493;
wire [15:0] slice_586;
wire [16:0] mulnw_5249;
wire [25:0] lsl_1342;
wire [47:0] addW_6005;
wire [17:0] slice_2098;
wire [7:0] slice_6761;
wire [17:0] slice_2854;
wire [15:0] slice_7517;
wire [98:0] concat_3610;
wire [66:0] concat_4366;
wire [32:0] lsl_459;
wire [34:0] addW_5122;
wire [66:0] concat_1215;
wire [39:0] mul_5878;
wire [17:0] slice_1971;
wire [7:0] slice_6634;
wire [32:0] slice_2727;
wire [64:0] slice_7390;
wire [13:0] slice_3483;
wire [33:0] add_4239;
wire [27:0] mul_332;
wire [7:0] slice_4995;
wire [31:0] slice_1088;
wire [41:0] subW_5751;
wire [15:0] mul_1844;
wire [39:0] mul_6507;
wire [15:0] slice_2600;
wire [15:0] mul_7263;
wire [17:0] slice_3356;
wire [17:0] add_4112;
wire [67:0] subW_205;
wire [7:0] slice_4868;
wire [31:0] slice_961;
wire [16:0] mulnw_5624;
wire [7:0] slice_1717;
wire [66:0] concat_6380;
wire [15:0] slice_2473;
wire [47:0] addW_7136;
wire [15:0] mul_3229;
wire [17:0] slice_3985;
wire [33:0] addW_78;
wire [71:0] subW_4741;
wire [16:0] mulnw_5497;
wire [7:0] slice_1590;
wire [31:0] slice_6253;
wire [15:0] slice_2346;
wire [134:0] subW_7009;
wire [7:0] slice_3102;
wire [13:0] slice_3858;
wire [16:0] slice_4614;
wire [15:0] slice_707;
wire [17:0] slice_5370;
wire [98:0] concat_1463;
wire [45:0] concat_6126;
wire [34:0] addW_2219;
wire [7:0] slice_6882;
wire [25:0] lsl_2975;
wire [13:0] slice_3731;
wire [63:0] slice_4487;
wire [32:0] slice_580;
wire [7:0] slice_5243;
wire [32:0] lsl_1336;
wire [45:0] concat_5999;
wire [31:0] slice_2092;
wire [7:0] slice_6755;
wire [19:0] addW_2848;
wire [25:0] lsl_7511;
wire [40:0] subW_3604;
wire [15:0] mul_4360;
wire [15:0] mul_453;
wire [17:0] slice_5116;
wire [15:0] mul_1209;
wire [17:0] slice_5872;
wire [19:0] addW_1965;
wire [26:0] add_6628;
wire [98:0] addW_2721;
wire [69:0] concat_7384;
wire [40:0] subW_3477;
wire [7:0] slice_4233;
wire [17:0] slice_326;
wire [26:0] add_4989;
wire [34:0] addW_1082;
wire [17:0] slice_5745;
wire [7:0] slice_1838;
wire [17:0] slice_6501;
wire [33:0] addW_2594;
wire [7:0] slice_7257;
wire [19:0] addW_3350;
wire [16:0] mulnw_4106;
wire [26:0] add_199;
wire [26:0] add_4862;
wire [31:0] slice_955;
wire [15:0] slice_5618;
wire [8:0] slice_1711;
wire [15:0] mul_6374;
wire [66:0] concat_2467;
wire [45:0] concat_7130;
wire [7:0] slice_3223;
wire [19:0] addW_3979;
wire [40:0] subW_4735;
wire [34:0] addW_828;
wire [33:0] add_5491;
wire [15:0] slice_1584;
wire [67:0] subW_6247;
wire [16:0] slice_2340;
wire [69:0] concat_7003;
wire [8:0] slice_3096;
wire [50:0] addW_3852;
wire [47:0] addW_4608;
wire [33:0] addW_701;
wire [31:0] slice_5364;
wire [40:0] subW_1457;
wire [13:0] slice_6120;
wire [41:0] subW_2213;
wire [26:0] add_6876;
wire [32:0] lsl_2969;
wire [130:0] concat_3725;
wire [134:0] subW_4481;
wire [129:0] addW_574;
wire [15:0] slice_5237;
wire [15:0] mul_1330;
wire [13:0] slice_5993;
wire [41:0] subW_2086;
wire [16:0] mulnw_6749;
wire [27:0] mul_2842;
wire [32:0] lsl_7505;
wire [35:0] mul_3598;
wire [7:0] slice_4354;
wire [7:0] slice_447;
wire [19:0] addW_5110;
wire [7:0] slice_1203;
wire [34:0] addW_5866;
wire [31:0] mul_1959;
wire [15:0] mulnw_6622;
wire [34:0] addW_2715;
wire [19:0] addW_7378;
wire [35:0] mul_3471;
wire [7:0] slice_4227;
wire [19:0] addW_320;
wire [15:0] mulnw_4983;
wire [15:0] mulnw_1076;
wire [31:0] slice_5739;
wire [15:0] slice_1832;
wire [34:0] addW_6495;
wire [41:0] subW_2588;
wire [26:0] add_7251;
wire [31:0] mul_3344;
wire [25:0] lsl_4100;
wire [16:0] mulnw_193;
wire [15:0] mulnw_4856;
wire [50:0] addW_949;
wire [130:0] addW_5612;
wire [33:0] mul_1705;
wire [7:0] slice_6368;
wire [15:0] mul_2461;
wire [13:0] slice_7124;
wire [15:0] slice_3217;
wire [31:0] mul_3973;
wire [41:0] subW_66;
wire [35:0] mul_4729;
wire [15:0] mulnw_822;
wire [7:0] slice_5485;
wire [32:0] slice_1578;
wire [26:0] add_6241;
wire [71:0] subW_2334;
wire [19:0] addW_6997;
wire [33:0] mul_3090;
wire [17:0] add_3846;
wire [45:0] concat_4602;
wire [41:0] subW_695;
wire [39:0] mul_5358;
wire [35:0] mul_1451;
wire [50:0] addW_6114;
wire [17:0] slice_2207;
wire [15:0] mulnw_6870;
wire [15:0] mul_2963;
wire [15:0] slice_3719;
wire [69:0] concat_4475;
wire [63:0] slice_568;
wire [32:0] slice_5231;
wire [7:0] slice_1324;
wire [130:0] concat_5987;
wire [17:0] slice_2080;
wire [7:0] slice_6743;
wire [17:0] slice_2836;
wire [15:0] mul_7499;
wire [13:0] slice_3592;
wire [26:0] add_4348;
wire [15:0] slice_441;
wire [27:0] mul_5104;
wire [26:0] add_1197;
wire [34:0] addW_5860;
wire [32:0] slice_1953;
wire [49:0] concat_6616;
wire [15:0] mulnw_2709;
wire [17:0] slice_7372;
wire [63:0] slice_3465;
wire [16:0] mulnw_4221;
wire [27:0] mul_314;
wire [49:0] concat_4977;
wire [8:0] slice_1070;
wire [34:0] addW_5733;
wire [33:0] addW_1826;
wire [41:0] subW_6489;
wire [17:0] slice_2582;
wire [15:0] mulnw_7245;
wire [32:0] slice_3338;
wire [32:0] lsl_4094;
wire [33:0] add_187;
wire [49:0] concat_4850;
wire [17:0] add_943;
wire [127:0] slice_5606;
wire [16:0] slice_1699;
wire [26:0] add_6362;
wire [7:0] slice_2455;
wire [47:0] addW_7118;
wire [33:0] addW_3211;
wire [31:0] slice_3967;
wire [17:0] slice_60;
wire [15:0] slice_4723;
wire [8:0] slice_816;
wire [8:0] slice_5479;
wire [63:0] slice_1572;
wire [16:0] mulnw_6235;
wire [40:0] subW_2328;
wire [17:0] slice_6991;
wire [32:0] slice_3084;
wire [16:0] mulnw_3840;
wire [13:0] slice_4596;
wire [17:0] slice_689;
wire [17:0] slice_5352;
wire [13:0] slice_1445;
wire [17:0] add_6108;
wire [31:0] slice_2201;
wire [49:0] concat_6864;
wire [7:0] slice_2957;
wire [25:0] lsl_3713;
wire [19:0] addW_4469;
wire [99:0] addW_562;
wire [98:0] addW_5225;
wire [15:0] slice_1318;
wire [15:0] slice_5981;
wire [31:0] slice_2074;
wire [15:0] slice_6737;
wire [19:0] addW_2830;
wire [7:0] slice_7493;
wire [33:0] add_3586;
wire [15:0] mulnw_4342;
wire [33:0] addW_435;
wire [15:0] slice_5098;
wire [15:0] mulnw_1191;
wire [15:0] mulnw_5854;
wire [26:0] add_1947;
wire [16:0] slice_6610;
wire [8:0] slice_2703;
wire [98:0] concat_7366;
wire [98:0] addW_3459;
wire [7:0] slice_4215;
wire [31:0] slice_308;
wire [16:0] slice_4971;
wire [17:0] add_1064;
wire [15:0] mulnw_5727;
wire [17:0] slice_1820;
wire [17:0] slice_6483;
wire [31:0] slice_2576;
wire [49:0] concat_7239;
wire [26:0] add_3332;
wire [31:0] mul_4088;
wire [7:0] slice_181;
wire [16:0] slice_4844;
wire [16:0] mulnw_937;
wire [131:0] concat_5600;
wire [15:0] mulnw_6356;
wire [26:0] add_2449;
wire [45:0] concat_7112;
wire [17:0] slice_3205;
wire [39:0] mul_3961;
wire [31:0] slice_54;
wire [47:0] addW_4717;
wire [17:0] add_810;
wire [33:0] mul_5473;
wire [66:0] concat_1566;
wire [33:0] add_6229;
wire [35:0] mul_2322;
wire [99:0] concat_6985;
wire [63:0] slice_3078;
wire [25:0] lsl_3834;
wire [47:0] addW_4590;
wire [31:0] slice_683;
wire [127:0] slice_5346;
wire [33:0] add_1439;
wire [16:0] mulnw_6102;
wire [34:0] addW_2195;
wire [16:0] slice_6858;
wire [15:0] slice_2951;
wire [32:0] lsl_3707;
wire [17:0] slice_4463;
wire [41:0] subW_556;
wire [34:0] addW_5219;
wire [32:0] slice_1312;
wire [25:0] lsl_5975;
wire [31:0] slice_2068;
wire [258:0] addW_6731;
wire [27:0] mul_2824;
wire [15:0] slice_7487;
wire [7:0] slice_3580;
wire [49:0] concat_4336;
wire [17:0] slice_429;
wire [25:0] lsl_5092;
wire [49:0] concat_1185;
wire [8:0] slice_5848;
wire [16:0] mulnw_1941;
wire [195:0] concat_6604;
wire [17:0] add_2697;
wire [40:0] subW_7360;
wire [34:0] addW_3453;
wire [15:0] slice_4209;
wire [133:0] subW_302;
wire [50:0] addW_4965;
wire [16:0] mulnw_1058;
wire [8:0] slice_5721;
wire [19:0] addW_1814;
wire [31:0] slice_6477;
wire [41:0] subW_2570;
wire [16:0] slice_7233;
wire [16:0] mulnw_3326;
wire [66:0] addW_4082;
wire [8:0] slice_175;
wire [131:0] concat_4838;
wire [25:0] lsl_931;
wire [17:0] slice_5594;
wire [262:0] subW_1687;
wire [49:0] concat_6350;
wire [15:0] mulnw_2443;
wire [13:0] slice_7106;
wire [19:0] addW_3199;
wire [17:0] slice_3955;
wire [41:0] subW_48;
wire [45:0] concat_4711;
wire [16:0] mulnw_804;
wire [31:0] slice_5467;
wire [15:0] mul_1560;
wire [7:0] slice_6223;
wire [15:0] slice_2316;
wire [33:0] add_6979;
wire [99:0] addW_3072;
wire [32:0] lsl_3828;
wire [45:0] concat_4584;
wire [41:0] subW_677;
wire [63:0] slice_5340;
wire [7:0] slice_1433;
wire [25:0] lsl_6096;
wire [15:0] mulnw_2189;
wire [65:0] concat_6852;
wire [33:0] addW_2945;
wire [15:0] mul_3701;
wire [99:0] concat_4457;
wire [17:0] slice_550;
wire [15:0] mulnw_5213;
wire [63:0] slice_1306;
wire [32:0] lsl_5969;
wire [50:0] addW_2062;
wire [31:0] slice_2818;
wire [32:0] slice_7481;
wire [7:0] slice_3574;
wire [16:0] slice_4330;
wire [19:0] addW_423;
wire [32:0] lsl_5086;
wire [16:0] slice_1179;
wire [17:0] add_5842;
wire [33:0] add_1935;
wire [67:0] subW_6598;
wire [16:0] mulnw_2691;
wire [35:0] mul_7354;
wire [15:0] mulnw_3447;
wire [257:0] addW_4203;
wire [70:0] subW_296;
wire [17:0] add_4959;
wire [15:0] slice_1052;
wire [17:0] add_5715;
wire [27:0] mul_1808;
wire [34:0] addW_6471;
wire [17:0] slice_2564;
wire [50:0] addW_7227;
wire [33:0] add_3320;
wire [130:0] concat_4076;
wire [33:0] mul_169;
wire [17:0] slice_4832;
wire [32:0] lsl_925;
wire [19:0] addW_5588;
wire [134:0] subW_1681;
wire [16:0] slice_6344;
wire [49:0] concat_2437;
wire [131:0] concat_7100;
wire [27:0] mul_3193;
wire [31:0] slice_3949;
wire [13:0] slice_4705;
wire [15:0] slice_798;
wire [39:0] mul_5461;
wire [7:0] slice_1554;
wire [8:0] slice_6217;
wire [47:0] addW_2310;
wire [7:0] slice_6973;
wire [41:0] subW_3066;
wire [31:0] mul_3822;
wire [13:0] slice_4578;
wire [17:0] slice_671;
wire [100:0] addW_5334;
wire [7:0] slice_1427;
wire [32:0] lsl_6090;
wire [8:0] slice_2183;
wire [19:0] addW_6846;
wire [17:0] slice_2939;
wire [511:0] slice_7602;
wire [7:0] slice_3695;
wire [33:0] add_4451;
wire [34:0] addW_544;
wire [8:0] slice_5207;
wire [66:0] concat_1300;
wire [15:0] mul_5963;
wire [17:0] add_2056;
wire [388:0] addW_6719;
wire [133:0] subW_2812;
wire [64:0] slice_7475;
wire [16:0] mulnw_3568;
wire [65:0] concat_4324;
wire [27:0] mul_417;
wire [15:0] mul_5080;
wire [65:0] concat_1173;
wire [16:0] mulnw_5836;
wire [7:0] slice_1929;
wire [26:0] add_6592;
wire [15:0] slice_2685;
wire [13:0] slice_7348;
wire [8:0] slice_3441;
wire [772:0] concat_4197;
wire [39:0] mul_290;
wire [16:0] mulnw_4953;
wire [16:0] slice_1046;
wire [16:0] mulnw_5709;
wire [17:0] slice_1802;
wire [15:0] mulnw_6465;
wire [31:0] slice_2558;
wire [17:0] add_7221;
wire [7:0] slice_3314;
wire [15:0] slice_4070;
wire [31:0] slice_163;
wire [19:0] addW_4826;
wire [31:0] mul_919;
wire [31:0] mul_5582;
wire [69:0] concat_1675;
wire [194:0] concat_6338;
wire [16:0] slice_2431;
wire [17:0] slice_7094;
wire [17:0] slice_3187;
wire [26:0] add_3943;
wire [17:0] slice_36;
wire [50:0] addW_4699;
wire [32:0] slice_792;
wire [17:0] slice_5455;
wire [26:0] add_1548;
wire [33:0] mul_6211;
wire [45:0] concat_2304;
wire [7:0] slice_6967;
wire [17:0] slice_3060;
wire [65:0] addW_3816;
wire [130:0] concat_4572;
wire [31:0] slice_665;
wire [41:0] subW_5328;
wire [16:0] mulnw_1421;
wire [31:0] mul_6084;
wire [17:0] add_2177;
wire [17:0] slice_6840;
wire [19:0] addW_2933;
wire [774:0] addW_7596;
wire [15:0] slice_3689;
wire [7:0] slice_4445;
wire [17:0] slice_538;
wire [17:0] add_5201;
wire [15:0] mul_1294;
wire [7:0] slice_5957;
wire [16:0] mulnw_2050;
wire [135:0] subW_6713;
wire [70:0] subW_2806;
wire [69:0] concat_7469;
wire [7:0] slice_3562;
wire [19:0] addW_4318;
wire [17:0] slice_411;
wire [7:0] slice_5074;
wire [19:0] addW_1167;
wire [15:0] slice_5830;
wire [8:0] slice_1923;
wire [16:0] mulnw_6586;
wire [33:0] addW_2679;
wire [33:0] add_7342;
wire [17:0] add_3435;
wire [261:0] subW_4191;
wire [17:0] slice_284;
wire [25:0] lsl_4947;
wire [31:0] slice_1040;
wire [15:0] slice_5703;
wire [19:0] addW_1796;
wire [8:0] slice_6459;
wire [31:0] slice_2552;
wire [16:0] mulnw_7215;
wire [8:0] slice_3308;
wire [25:0] lsl_4064;
wire [39:0] mul_157;
wire [31:0] mul_4820;
wire [16:0] slice_913;
wire [31:0] slice_5576;
wire [19:0] addW_1669;
wire [67:0] subW_6332;
wire [19:0] addW_7088;
wire [19:0] addW_3181;
wire [16:0] mulnw_3937;
wire [63:0] slice_30;
wire [17:0] add_4693;
wire [26:0] add_786;
wire [31:0] slice_5449;
wire [15:0] mulnw_1542;
wire [31:0] slice_6205;
wire [13:0] slice_2298;
wire [16:0] mulnw_6961;
wire [34:0] addW_3054;
wire [130:0] concat_3810;
wire [15:0] slice_4566;
wire [31:0] slice_659;
wire [17:0] slice_5322;
wire [7:0] slice_1415;
wire [65:0] addW_6078;
wire [16:0] mulnw_2171;
wire [65:0] concat_6834;
wire [27:0] mul_2927;
wire [264:0] subW_7590;
wire [33:0] addW_3683;
wire [7:0] slice_4439;
wire [19:0] addW_532;
wire [16:0] mulnw_5195;
wire [7:0] slice_1288;
wire [15:0] slice_5951;
wire [25:0] lsl_2044;
wire [70:0] subW_6707;
wire [39:0] mul_2800;
wire [19:0] addW_7463;
wire [15:0] slice_3556;
wire [17:0] slice_4312;
wire [19:0] addW_405;
wire [15:0] slice_5068;
wire [17:0] slice_1161;
wire [32:0] slice_5824;
wire [33:0] mul_1917;
wire [33:0] add_6580;
wire [41:0] subW_2673;
wire [7:0] slice_7336;
wire [16:0] mulnw_3429;
wire [133:0] concat_4185;
wire [34:0] addW_278;
wire [32:0] lsl_4941;
wire [50:0] addW_1034;
wire [16:0] slice_5697;
wire [27:0] mul_1790;
wire [17:0] add_6453;
wire [255:0] slice_2546;
wire [25:0] lsl_7209;
wire [33:0] mul_3302;
wire [32:0] lsl_4058;
wire [17:0] slice_151;
wire [31:0] slice_4814;
wire [47:0] addW_907;
wire [39:0] mul_5570;
wire [17:0] slice_1663;
wire [26:0] add_6326;
wire [71:0] subW_2419;
wire [31:0] mul_7082;
wire [27:0] mul_3175;
wire [33:0] add_3931;
wire [16:0] mulnw_4687;
wire [16:0] mulnw_780;
wire [39:0] mul_5443;
wire [49:0] concat_1536;
wire [39:0] mul_6199;
wire [50:0] addW_2292;
wire [7:0] slice_6955;
wire [17:0] slice_3048;
wire [15:0] slice_3804;
wire [25:0] lsl_4560;
wire [51:0] addW_653;
wire [34:0] addW_5316;
wire [15:0] slice_1409;
wire [130:0] concat_6072;
wire [15:0] slice_2165;
wire [19:0] addW_6828;
wire [17:0] slice_2921;
wire [134:0] subW_7584;
wire [17:0] slice_3677;
wire [16:0] mulnw_4433;
wire [27:0] mul_526;
wire [15:0] slice_5189;
wire [26:0] add_1282;
wire [33:0] addW_5945;
wire [32:0] lsl_2038;
wire [39:0] mul_6701;
wire [17:0] slice_2794;
wire [17:0] slice_7457;
wire [32:0] slice_3550;
wire [65:0] concat_4306;
wire [27:0] mul_399;
wire [32:0] slice_5062;
wire [65:0] concat_1155;
wire [26:0] add_5818;
wire [15:0] slice_1911;
wire [7:0] slice_6574;
wire [17:0] slice_2667;
wire [7:0] slice_7330;
wire [15:0] slice_3423;
wire [17:0] slice_4179;
wire [17:0] slice_272;
wire [31:0] mul_4935;
wire [17:0] add_1028;
wire [71:0] subW_5691;
wire [63:0] slice_1784;
wire [16:0] mulnw_6447;
wire [389:0] addW_2540;
wire [32:0] lsl_7203;
wire [15:0] slice_3296;
wire [15:0] mul_4052;
wire [31:0] slice_145;
wire [39:0] mul_4808;
wire [45:0] concat_901;
wire [17:0] slice_5564;
wire [99:0] concat_1657;
wire [16:0] mulnw_6320;
wire [40:0] subW_2413;
wire [31:0] slice_7076;
wire [63:0] slice_3169;
wire [7:0] slice_3925;
wire [25:0] lsl_4681;
wire [33:0] add_774;
wire [17:0] slice_5437;
wire [16:0] slice_1530;
wire [17:0] slice_6193;
wire [17:0] add_2286;
wire [15:0] slice_6949;
wire [19:0] addW_3042;
wire [25:0] lsl_3798;
wire [32:0] lsl_4554;
wire [49:0] concat_647;
wire [15:0] slice_5310;
wire [16:0] slice_1403;
wire [15:0] slice_6066;
wire [16:0] slice_2159;
wire [17:0] slice_6822;
wire [19:0] addW_2915;
wire [69:0] concat_7578;
wire [19:0] addW_3671;
wire [7:0] slice_4427;
wire [15:0] slice_520;
wire [33:0] addW_5183;
wire [15:0] mulnw_1276;
wire [17:0] slice_5939;
wire [31:0] mul_2032;
wire [17:0] slice_6695;
wire [34:0] addW_2788;
wire [98:0] concat_7451;
wire [98:0] addW_3544;
wire [19:0] addW_4300;
wire [63:0] slice_393;
wire [32:0] slice_5056;
wire [19:0] addW_1149;
wire [16:0] mulnw_5812;
wire [25:0] lsl_1905;
wire [8:0] slice_6568;
wire [31:0] slice_2661;
wire [16:0] mulnw_7324;
wire [33:0] addW_3417;
wire [19:0] addW_4173;
wire [19:0] addW_266;
wire [66:0] addW_4929;
wire [16:0] mulnw_1022;
wire [40:0] subW_5685;
wire [69:0] concat_1778;
wire [15:0] slice_6441;
wire [135:0] subW_2534;
wire [31:0] mul_7197;
wire [25:0] lsl_3290;
wire [7:0] slice_4046;
wire [39:0] mul_139;
wire [17:0] slice_4802;
wire [13:0] slice_895;
wire [31:0] slice_5558;
wire [33:0] add_1651;
wire [33:0] add_6314;
wire [35:0] mul_2407;
wire [39:0] mul_7070;
wire [69:0] concat_3163;
wire [8:0] slice_3919;
wire [32:0] lsl_4675;
wire [7:0] slice_768;
wire [13:0] slice_5431;
wire [65:0] concat_1524;
wire [31:0] slice_6187;
wire [16:0] mulnw_2280;
wire [66:0] concat_6943;
wire [27:0] mul_3036;
wire [32:0] lsl_3792;
wire [15:0] mul_4548;
wire [15:0] slice_641;
wire [25:0] lsl_5304;
wire [259:0] concat_1397;
wire [25:0] lsl_6060;
wire [31:0] slice_2153;
wire [31:0] slice_6816;
wire [27:0] mul_2909;
wire [19:0] addW_7572;
wire [27:0] mul_3665;
wire [15:0] slice_4421;
wire [25:0] lsl_514;
wire [41:0] subW_5177;
wire [49:0] concat_1270;
wire [19:0] addW_5933;
wire [16:0] slice_2026;
wire [34:0] addW_6689;
wire [41:0] subW_2782;
wire [40:0] subW_7445;
wire [34:0] addW_3538;
wire [17:0] slice_4294;
wire [66:0] concat_387;
wire [17:0] slice_1143;
wire [33:0] add_5806;
wire [32:0] lsl_1899;
wire [33:0] mul_6562;
wire [41:0] subW_2655;
wire [7:0] slice_7318;
wire [41:0] subW_3411;
wire [31:0] mul_4167;
wire [27:0] mul_260;
wire [131:0] concat_4923;
wire [25:0] lsl_1016;
wire [35:0] mul_5679;
wire [19:0] addW_1772;
wire [129:0] addW_6435;
wire [70:0] subW_2528;
wire [66:0] addW_7191;
wire [32:0] lsl_3284;
wire [15:0] slice_4040;
wire [17:0] slice_133;
wire [31:0] slice_4796;
wire [47:0] addW_889;
wire [26:0] add_5552;
wire [7:0] slice_1645;
wire [7:0] slice_6308;
wire [15:0] slice_2401;
wire [17:0] slice_7064;
wire [19:0] addW_3157;
wire [33:0] mul_3913;
wire [31:0] mul_4669;
wire [8:0] slice_762;
wire [68:0] subW_5425;
wire [19:0] addW_1518;
wire [39:0] mul_6181;
wire [25:0] lsl_2274;
wire [15:0] mul_6937;
wire [15:0] slice_3030;
wire [15:0] mul_3786;
wire [7:0] slice_4542;
wire [65:0] concat_635;
wire [32:0] lsl_5298;
wire [31:0] slice_1391;
wire [32:0] lsl_6054;
wire [50:0] addW_2147;
wire [70:0] subW_6810;
wire [63:0] slice_2903;
wire [17:0] slice_7566;
wire [17:0] slice_3659;
wire [66:0] concat_4415;
wire [32:0] lsl_508;
wire [17:0] slice_5171;
wire [16:0] slice_1264;
wire [27:0] mul_5927;
wire [47:0] addW_2020;
wire [34:0] addW_6683;
wire [17:0] slice_2776;
wire [35:0] mul_7439;
wire [15:0] mulnw_3532;
wire [31:0] slice_4288;
wire [15:0] mul_381;
wire [519:0] subW_5044;
wire [13:0] slice_1137;
wire [7:0] slice_5800;
wire [15:0] mul_1893;
wire [31:0] slice_6556;
wire [17:0] slice_2649;
wire [15:0] slice_7312;
wire [17:0] slice_3405;
wire [32:0] slice_4161;
wire [15:0] slice_254;
wire [17:0] slice_4917;
wire [32:0] lsl_1010;
wire [15:0] slice_5673;
wire [17:0] slice_1766;
wire [127:0] slice_6429;
wire [39:0] mul_2522;
wire [130:0] concat_7185;
wire [15:0] mul_3278;
wire [33:0] addW_4034;
wire [13:0] slice_127;
wire [26:0] add_4790;
wire [45:0] concat_883;
wire [16:0] mulnw_5546;
wire [7:0] slice_1639;
wire [8:0] slice_6302;
wire [47:0] addW_2395;
wire [31:0] slice_7058;
wire [17:0] slice_3151;
wire [32:0] slice_3907;
assign addW_4663 = slice_4576 + slice_4491;
assign mul_756 = slice_752 * slice_755;
assign add_5419 = lsl_5410 + add_5418;
assign slice_1512 = slice_1507[17:0];
assign slice_6175 = slice_6171[17:0];
assign lsl_2268 = mulnw_2267 << 16;
assign slice_6931 = slice_6909[7:0];
assign lsl_3024 = add_3023 << 8;
assign slice_3780 = slice_3767[7:0];
assign slice_4536 = mul_4535[31:16];
assign addW_629 = slice_624 + slice_621;
assign mul_5292 = slice_5286 * slice_5288;
assign addW_1385 = concat_1379 + subW_1384;
assign mul_6048 = slice_6042 * slice_6044;
assign add_2141 = mulnw_2138 + mulnw_2140;
assign mul_6804 = addW_6802 * addW_6803;
assign concat_2897 = {addW_2895,slice_2896};
assign concat_7560 = {concat_7518,slice_7559};
assign addW_3653 = slice_3648 + slice_3642;
assign mul_4409 = slice_4403 * slice_4405;
assign mul_502 = slice_496 * slice_498;
assign slice_5165 = slice_5146[31:0];
assign concat_1258 = {addW_1256,slice_1257};
assign slice_5921 = mul_5912[17:0];
assign concat_2014 = {mul_2009,slice_2013};
assign mulnw_6677 = slice_6670 * slice_6676;
assign slice_2770 = addW_2729[31:0];
assign slice_7433 = slice_7432[31:18];
assign slice_3526 = slice_3505[16:8];
assign subW_4282 = concat_4281 - concat_4243;
assign slice_375 = slice_353[7:0];
assign subW_5038 = concat_5037 - concat_4485;
assign addW_1131 = concat_1043 + subW_1130;
assign slice_5794 = slice_5784[16:8];
assign slice_1887 = slice_1873[7:0];
assign mul_6550 = addW_6548 * addW_6549;
assign slice_2643 = slice_2642[63:32];
assign slice_7306 = slice_7305[32:16];
assign slice_3399 = slice_3380[31:0];
assign add_4155 = lsl_4153 + mul_4154;
assign lsl_248 = add_247 << 8;
assign addW_4911 = slice_4906 + slice_4902;
assign mul_1004 = slice_1002 * slice_1003;
assign addW_5667 = concat_5661 + subW_5666;
assign concat_1760 = {concat_1740,slice_1759};
assign concat_6423 = {addW_6421,slice_6422};
assign slice_2516 = addW_2512[17:0];
assign slice_7179 = mul_7148[15:0];
assign slice_3272 = slice_3258[7:0];
assign slice_4028 = mul_4019[17:0];
assign subW_121 = subW_120 - concat_69;
assign mulnw_4784 = slice_4783 * slice_4780;
assign slice_877 = slice_876[31:18];
assign add_5540 = lsl_5531 + add_5539;
assign mulnw_1633 = slice_1626 * slice_1632;
assign mul_6296 = slice_6293 * slice_6295;
assign concat_2389 = {mul_2384,slice_2388};
assign add_7052 = lsl_7050 + mul_7051;
assign concat_3145 = {concat_3125,slice_3144};
assign slice_3901 = concat_3810[63:0];
assign concat_4657 = {addW_4655,slice_4656};
assign addW_750 = slice_661 + slice_575;
assign slice_5413 = slice_5387[7:0];
assign concat_1506 = {addW_1504,slice_1505};
assign slice_6169 = slice_5904[127:0];
assign mul_2262 = slice_2260 * slice_2261;
assign add_6925 = lsl_6923 + mul_6924;
assign lsl_3018 = mulnw_3017 << 16;
assign slice_3774 = mul_3773[31:16];
assign addW_4530 = slice_4510 + slice_4492;
assign slice_623 = slice_618[17:0];
assign slice_5286 = slice_5273[7:0];
assign concat_1379 = {mul_1374,slice_1378};
assign slice_6042 = slice_6029[7:0];
assign mulnw_2135 = slice_2133 * slice_2134;
assign slice_6798 = addW_6794[17:0];
assign mul_2891 = slice_2885 * slice_2887;
assign add_7554 = lsl_7545 + add_7553;
assign mul_3647 = slice_3642 * slice_3646;
assign slice_4403 = slice_4381[7:0];
assign slice_496 = slice_482[7:0];
assign subW_5159 = subW_5158 - mul_5152;
assign addW_1252 = slice_1247 + slice_1244;
assign addW_5915 = slice_5910 + slice_5903;
assign slice_2008 = slice_2007[31:18];
assign slice_6671 = slice_6650[16:8];
assign addW_2764 = add_2750 + add_2763;
assign add_7427 = lsl_7418 + add_7426;
assign add_3520 = mulnw_3517 + mulnw_3519;
assign mul_4276 = addW_4274 * addW_4275;
assign add_369 = lsl_367 + mul_368;
assign concat_5032 = {addW_5030,slice_5031};
assign subW_1125 = subW_1124 - concat_1103;
assign mul_5788 = slice_5784 * slice_5787;
assign slice_1881 = mul_1880[31:16];
assign slice_6544 = slice_6540[17:0];
assign slice_2637 = concat_2591[31:0];
assign slice_7300 = concat_7299[257:129];
assign subW_3393 = subW_3392 - mul_3386;
assign mulnw_4149 = slice_4148 * slice_4145;
assign lsl_242 = mulnw_241 << 16;
assign mul_4905 = slice_4902 * slice_4904;
assign slice_998 = addW_997[32:16];
assign concat_5661 = {mul_5656,slice_5660};
assign subW_1754 = mul_1753 - mul_1745;
assign slice_6417 = mul_6408[17:0];
assign addW_2510 = slice_2468 + slice_2427;
assign lsl_7173 = add_7172 << 8;
assign slice_3266 = mul_3265[31:16];
assign addW_4022 = slice_4017 + slice_4013;
assign add_115 = lsl_106 + add_114;
assign add_4778 = lsl_4769 + add_4777;
assign slice_871 = slice_870[63:32];
assign slice_5534 = slice_5524[7:0];
assign slice_1627 = slice_1622[15:8];
assign slice_6290 = concat_6289[63:32];
assign slice_2383 = slice_2382[31:18];
assign mulnw_7046 = slice_7045 * slice_7042;
assign subW_3139 = mul_3138 - mul_3130;
assign addW_3895 = concat_3874 + subW_3894;
assign slice_4651 = mul_4620[15:0];
assign slice_744 = concat_698[31:0];
assign slice_5407 = slice_5389[15:8];
assign addW_1500 = slice_1495 + slice_1492;
assign slice_6163 = concat_6072[63:0];
assign slice_2256 = addW_2255[129:65];
assign mulnw_6919 = slice_6918 * slice_6915;
assign mul_3012 = slice_3006 * slice_3008;
assign addW_3768 = slice_3748 + slice_3730;
assign slice_4524 = mul_4515[17:0];
assign concat_617 = {addW_615,slice_616};
assign slice_5280 = mul_5279[31:16];
assign slice_1373 = addW_1372[33:18];
assign slice_6036 = mul_6035[31:16];
assign lsl_2129 = add_2128 << 8;
assign addW_6792 = slice_6772 + slice_6729;
assign slice_2885 = slice_2863[7:0];
assign slice_7548 = slice_7522[7:0];
assign slice_3641 = slice_3640[63:32];
assign add_4397 = lsl_4395 + mul_4396;
assign slice_490 = mul_489[31:16];
assign slice_5153 = mul_5152[35:18];
assign slice_1246 = slice_1241[17:0];
assign mul_5909 = slice_5903 * slice_5908;
assign addW_2002 = concat_1996 + subW_2001;
assign add_6665 = mulnw_6662 + mulnw_6664;
assign mulnw_2758 = slice_2751 * slice_2757;
assign slice_7421 = slice_7395[7:0];
assign mulnw_3514 = slice_3512 * slice_3513;
assign slice_4270 = addW_4266[17:0];
assign mulnw_363 = slice_362 * slice_359;
assign slice_5026 = mul_5017[17:0];
assign subW_1119 = mul_1118 - mul_1110;
assign addW_5782 = slice_5695 + slice_5609;
assign slice_1875 = addW_1874[65:33];
assign slice_6538 = slice_6518[31:0];
assign addW_2631 = concat_2603 + addW_2630;
assign concat_7294 = {addW_7292,slice_7293};
assign slice_3387 = mul_3386[35:18];
assign add_4143 = lsl_4134 + add_4142;
assign mul_236 = slice_230 * slice_232;
assign slice_4899 = concat_4898[63:32];
assign addW_992 = concat_986 + subW_991;
assign slice_5655 = slice_5654[31:18];
assign mul_1748 = slice_1746 * slice_1747;
assign addW_6411 = slice_6406 + slice_6402;
assign addW_2504 = add_2490 + add_2503;
assign lsl_7167 = mulnw_7166 << 16;
assign slice_3260 = addW_3259[65:33];
assign mul_4016 = slice_4013 * slice_4015;
assign slice_109 = slice_79[7:0];
assign slice_4772 = slice_4762[7:0];
assign addW_865 = concat_571 + subW_864;
assign slice_5528 = slice_5518[16:8];
assign slice_1621 = slice_1616[15:0];
assign mul_6284 = addW_6282 * addW_6283;
assign addW_2377 = concat_2349 + addW_2376;
assign add_7040 = lsl_7031 + add_7039;
assign mul_3133 = slice_3131 * slice_3132;
assign subW_3889 = subW_3888 - mul_3882;
assign lsl_4645 = add_4644 << 8;
assign addW_738 = concat_710 + addW_737;
assign mulnw_5401 = slice_5394 * slice_5400;
assign slice_1494 = slice_1488[17:0];
assign addW_6157 = concat_6136 + subW_6156;
assign concat_6913 = {mul_6908,slice_6912};
assign slice_3006 = slice_2992[7:0];
assign slice_3762 = mul_3753[17:0];
assign addW_4518 = slice_4513 + slice_4509;
assign mul_611 = slice_605 * slice_607;
assign slice_5274 = addW_5233[32:0];
assign concat_1367 = {addW_1365,slice_1366};
assign addW_6030 = slice_6010 + slice_5992;
assign lsl_2123 = mulnw_2122 << 16;
assign subW_6786 = subW_6785 - mul_6779;
assign add_2879 = lsl_2877 + mul_2878;
assign slice_7542 = slice_7524[15:8];
assign subW_3635 = subW_3634 - concat_3546;
assign mulnw_4391 = slice_4390 * slice_4387;
assign slice_484 = addW_483[64:32];
assign slice_5147 = slice_5146[63:32];
assign concat_1240 = {addW_1238,slice_1239};
assign slice_5903 = slice_5902[31:18];
assign concat_1996 = {mul_1991,slice_1995};
assign mulnw_6659 = slice_6657 * slice_6658;
assign slice_2752 = slice_2731[16:8];
assign slice_7415 = slice_7397[15:8];
assign slice_3508 = addW_3504[15:0];
assign addW_4264 = slice_4244 + slice_4201;
assign concat_357 = {mul_352,slice_356};
assign addW_5020 = slice_5015 + slice_5011;
assign mul_1113 = slice_1111 * slice_1112;
assign subW_5776 = subW_5775 - concat_5754;
assign slice_1869 = concat_1868[127:64];
assign mul_6532 = addW_6530 * addW_6531;
assign add_2625 = mulnw_2622 + mulnw_2624;
assign slice_7288 = mul_7279[17:0];
assign slice_3381 = slice_3380[63:32];
assign slice_4137 = slice_4127[7:0];
assign slice_230 = slice_216[7:0];
assign mul_4893 = addW_4891 * addW_4892;
assign concat_986 = {mul_981,slice_985};
assign addW_5649 = concat_5621 + addW_5648;
assign slice_1742 = slice_1741[31:18];
assign mul_6405 = slice_6402 * slice_6404;
assign mulnw_2498 = slice_2491 * slice_2497;
assign mul_7161 = slice_7155 * slice_7157;
assign slice_3254 = concat_3253[127:64];
assign slice_4010 = mul_4001[17:0];
assign slice_103 = slice_82[15:8];
assign slice_4766 = slice_4755[16:8];
assign subW_859 = subW_858 - concat_745;
assign mul_5522 = slice_5518 * slice_5521;
assign concat_1615 = {addW_1613,slice_1614};
assign slice_6278 = slice_6274[17:0];
assign add_2371 = mulnw_2368 + mulnw_2370;
assign slice_7034 = slice_7024[7:0];
assign slice_3127 = slice_3126[31:18];
assign slice_3883 = mul_3882[35:18];
assign lsl_4639 = mulnw_4638 << 16;
assign add_732 = mulnw_729 + mulnw_731;
assign slice_5395 = slice_5390[15:8];
assign slice_1488 = slice_1487[63:32];
assign subW_6151 = subW_6150 - mul_6144;
assign addW_2244 = concat_2156 + subW_2243;
assign slice_6907 = slice_6906[32:16];
assign slice_3000 = mul_2999[31:16];
assign addW_3756 = slice_3751 + slice_3747;
assign mul_4512 = slice_4509 * slice_4511;
assign slice_605 = slice_583[7:0];
assign addW_5268 = add_5254 + add_5267;
assign addW_1361 = slice_1356 + slice_1353;
assign slice_6024 = mul_6015[17:0];
assign mul_2117 = slice_2115 * slice_2116;
assign slice_6780 = mul_6779[35:18];
assign mulnw_2873 = slice_2872 * slice_2869;
assign mulnw_7536 = slice_7529 * slice_7535;
assign subW_3629 = concat_3628 - concat_3590;
assign concat_4385 = {mul_4380,slice_4384};
assign slice_478 = concat_477[127:64];
assign slice_5141 = concat_5117[31:0];
assign addW_1234 = slice_1229 + slice_1226;
assign slice_5897 = concat_5605[127:0];
assign slice_1990 = slice_1989[31:18];
assign slice_6653 = slice_6649[15:0];
assign add_2746 = mulnw_2743 + mulnw_2745;
assign mulnw_7409 = slice_7402 * slice_7408;
assign addW_3502 = slice_3482 + slice_3463;
assign subW_4258 = subW_4257 - mul_4251;
assign slice_351 = addW_350[32:16];
assign mul_5014 = slice_5011 * slice_5013;
assign slice_1107 = addW_1106[33:18];
assign subW_5770 = mul_5769 - mul_5761;
assign concat_1863 = {addW_1861,slice_1862};
assign slice_6526 = slice_6522[17:0];
assign mulnw_2619 = slice_2617 * slice_2618;
assign addW_7282 = slice_7277 + slice_7273;
assign slice_3375 = slice_3374[127:64];
assign slice_4131 = slice_4122[16:8];
assign slice_224 = mul_223[31:16];
assign slice_4887 = slice_4883[17:0];
assign slice_980 = slice_979[31:18];
assign add_5643 = mulnw_5640 + mulnw_5642;
assign add_1736 = lsl_1727 + add_1735;
assign slice_6399 = concat_6398[63:32];
assign slice_2492 = slice_2471[16:8];
assign slice_7155 = slice_7142[7:0];
assign concat_3248 = {addW_3246,slice_3247};
assign addW_4004 = slice_3999 + slice_3994;
assign mulnw_97 = slice_89 * slice_96;
assign mul_4760 = slice_4755 * slice_4759;
assign subW_853 = concat_852 - concat_791;
assign addW_5516 = slice_5429 + slice_5343;
assign mul_1609 = slice_1603 * slice_1605;
assign slice_6272 = slice_6252[31:0];
assign mulnw_2365 = slice_2363 * slice_2364;
assign slice_7028 = slice_7017[16:8];
assign add_3121 = lsl_3112 + add_3120;
assign addW_3877 = slice_3857 + slice_3817;
assign mul_4633 = slice_4627 * slice_4629;
assign mulnw_726 = slice_724 * slice_725;
assign slice_5389 = addW_5384[15:0];
assign subW_1482 = concat_1481 - concat_1443;
assign slice_6145 = mul_6144[35:18];
assign subW_2238 = subW_2237 - concat_2216;
assign concat_6901 = {concat_6814,slice_6900};
assign slice_2994 = addW_2993[64:32];
assign mul_3750 = slice_3747 * slice_3749;
assign slice_4506 = mul_4497[17:0];
assign add_599 = lsl_597 + mul_598;
assign mulnw_5262 = slice_5255 * slice_5261;
assign slice_1355 = slice_1350[17:0];
assign addW_6018 = slice_6013 + slice_6009;
assign slice_2111 = addW_2110[32:16];
assign slice_6774 = slice_6733[31:0];
assign concat_2867 = {mul_2862,slice_2866};
assign slice_7530 = slice_7525[15:8];
assign mul_3623 = addW_3621 * addW_3622;
assign slice_4379 = slice_4378[32:16];
assign concat_472 = {addW_470,slice_471};
assign addW_5135 = concat_5129 + subW_5134;
assign slice_1228 = slice_1222[17:0];
assign addW_5891 = concat_5781 + subW_5890;
assign slice_1984 = slice_1983[127:64];
assign slice_6647 = addW_6605[32:0];
assign mulnw_2740 = slice_2738 * slice_2739;
assign slice_7403 = slice_7398[15:8];
assign subW_3496 = subW_3495 - mul_3489;
assign slice_4252 = mul_4251[35:18];
assign concat_345 = {addW_343,slice_344};
assign slice_5008 = concat_5007[65:33];
assign addW_1101 = concat_1095 + subW_1100;
assign mul_5764 = slice_5762 * slice_5763;
assign mul_1857 = slice_1851 * slice_1853;
assign slice_6520 = slice_6519[31:18];
assign lsl_2613 = add_2612 << 8;
assign mul_7276 = slice_7273 * slice_7275;
assign subW_3369 = subW_3368 - concat_3079;
assign mul_4125 = slice_4122 * slice_4124;
assign slice_218 = addW_217[64:32];
assign slice_4881 = slice_4839[31:0];
assign addW_974 = concat_968 + subW_973;
assign mulnw_5637 = slice_5635 * slice_5636;
assign slice_1730 = slice_1704[7:0];
assign mul_6393 = addW_6391 * addW_6392;
assign add_2486 = mulnw_2483 + mulnw_2485;
assign slice_7149 = mul_7148[31:16];
assign mul_3242 = slice_3236 * slice_3238;
assign mul_3998 = slice_3994 * slice_3997;
assign mulnw_91 = slice_89 * slice_90;
assign slice_4754 = slice_4753[64:32];
assign mul_847 = addW_845 * addW_846;
assign subW_5510 = subW_5509 - concat_5466;
assign slice_1603 = slice_1581[7:0];
assign mul_6266 = addW_6264 * addW_6265;
assign lsl_2359 = add_2358 << 8;
assign mul_7022 = slice_7017 * slice_7021;
assign slice_3115 = slice_3089[7:0];
assign slice_3871 = mul_3862[17:0];
assign slice_4627 = slice_4614[7:0];
assign lsl_720 = add_719 << 8;
assign concat_5383 = {concat_5363,slice_5382};
assign mul_1476 = addW_1474 * addW_1475;
assign addW_6139 = slice_6119 + slice_6079;
assign subW_2232 = mul_2231 - mul_2223;
assign subW_6895 = concat_6894 - concat_6834;
assign slice_2988 = concat_2987[127:64];
assign slice_3744 = mul_3735[17:0];
assign addW_4500 = slice_4495 + slice_4489;
assign mulnw_593 = slice_592 * slice_589;
assign slice_5256 = slice_5235[16:8];
assign concat_1349 = {addW_1347,slice_1348};
assign mul_6012 = slice_6009 * slice_6011;
assign addW_2105 = concat_2099 + subW_2104;
assign addW_6768 = add_6754 + add_6767;
assign slice_2861 = addW_2860[32:16];
assign slice_7524 = slice_7519[15:0];
assign slice_3617 = addW_3613[17:0];
assign concat_4373 = {concat_4286,slice_4372};
assign mul_466 = slice_460 * slice_462;
assign concat_5129 = {mul_5124,slice_5128};
assign slice_1222 = slice_1221[63:32];
assign subW_5885 = subW_5884 - concat_5863;
assign subW_1978 = concat_1977 - concat_1783;
assign add_6641 = lsl_6639 + mul_6640;
assign slice_2734 = slice_2730[15:0];
assign slice_7397 = slice_7391[15:0];
assign slice_3490 = mul_3489[35:18];
assign slice_4246 = slice_4205[31:0];
assign addW_339 = slice_334 + slice_331;
assign add_5002 = lsl_5000 + mul_5001;
assign concat_1095 = {mul_1090,slice_1094};
assign slice_5758 = addW_5757[33:18];
assign slice_1851 = slice_1829[7:0];
assign subW_6514 = subW_6513 - concat_6492;
assign lsl_2607 = mulnw_2606 << 16;
assign slice_7270 = concat_7269[65:33];
assign subW_3363 = concat_3362 - concat_3168;
assign slice_4119 = mul_4088[15:0];
assign add_4875 = lsl_4873 + mul_4874;
assign concat_968 = {mul_963,slice_967};
assign lsl_5631 = add_5630 << 8;
assign slice_1724 = slice_1706[15:8];
assign slice_6387 = slice_6383[17:0];
assign mulnw_2480 = slice_2478 * slice_2479;
assign addW_7143 = slice_7123 + slice_7105;
assign slice_3236 = slice_3214[7:0];
assign slice_3992 = addW_3905[63:0];
assign slice_85 = mul_84[31:16];
assign slice_4748 = concat_4657[63:0];
assign slice_841 = addW_837[17:0];
assign add_5504 = lsl_5495 + add_5503;
assign add_1597 = lsl_1595 + mul_1596;
assign slice_6260 = slice_6256[17:0];
assign lsl_2353 = mulnw_2352 << 16;
assign slice_7016 = slice_7015[64:32];
assign slice_3109 = slice_3091[15:8];
assign addW_3865 = slice_3860 + slice_3856;
assign slice_4621 = mul_4620[31:16];
assign lsl_714 = mulnw_713 << 16;
assign subW_5377 = mul_5376 - mul_5368;
assign slice_1470 = addW_1466[17:0];
assign slice_6133 = mul_6124[17:0];
assign mul_2226 = slice_2224 * slice_2225;
assign add_6889 = lsl_6887 + mul_6888;
assign concat_2982 = {addW_2980,slice_2981};
assign addW_3738 = slice_3733 + slice_3728;
assign mul_4494 = slice_4489 * slice_4493;
assign concat_587 = {mul_582,slice_586};
assign add_5250 = mulnw_5247 + mulnw_5249;
assign mul_1343 = slice_1337 * slice_1339;
assign slice_6006 = mul_5997[17:0];
assign concat_2099 = {mul_2094,slice_2098};
assign mulnw_6762 = slice_6755 * slice_6761;
assign concat_2855 = {addW_2853,slice_2854};
assign concat_7518 = {addW_7516,slice_7517};
assign addW_3611 = slice_3591 + slice_3550;
assign subW_4367 = concat_4366 - concat_4306;
assign slice_460 = slice_438[7:0];
assign slice_5123 = addW_5122[33:18];
assign subW_1216 = concat_1215 - concat_1155;
assign subW_5879 = mul_5878 - mul_5870;
assign concat_1972 = {addW_1970,slice_1971};
assign mulnw_6635 = slice_6634 * slice_6631;
assign slice_2728 = slice_2727[32:16];
assign slice_7391 = slice_7390[64:32];
assign slice_3484 = slice_3465[31:0];
assign addW_4240 = add_4226 + add_4239;
assign slice_333 = slice_328[17:0];
assign mulnw_4996 = slice_4995 * slice_4992;
assign slice_1089 = slice_1088[31:18];
assign addW_5752 = concat_5746 + subW_5751;
assign add_1845 = lsl_1843 + mul_1844;
assign subW_6508 = mul_6507 - mul_6499;
assign mul_2601 = slice_2599 * slice_2600;
assign add_7264 = lsl_7262 + mul_7263;
assign concat_3357 = {addW_3355,slice_3356};
assign lsl_4113 = add_4112 << 8;
assign subW_206 = subW_205 - concat_162;
assign mulnw_4869 = slice_4868 * slice_4865;
assign slice_962 = slice_961[31:18];
assign lsl_5625 = mulnw_5624 << 16;
assign mulnw_1718 = slice_1711 * slice_1717;
assign slice_6381 = addW_6339[31:0];
assign slice_2474 = slice_2470[15:0];
assign slice_7137 = mul_7128[17:0];
assign add_3230 = lsl_3228 + mul_3229;
assign concat_3986 = {addW_3984,slice_3985};
assign slice_79 = addW_78[32:16];
assign addW_4742 = concat_4721 + subW_4741;
assign addW_835 = slice_792 + slice_751;
assign slice_5498 = slice_5472[7:0];
assign mulnw_1591 = slice_1590 * slice_1587;
assign slice_6254 = slice_6253[31:18];
assign mul_2347 = slice_2345 * slice_2346;
assign subW_7010 = subW_7009 - concat_6899;
assign mulnw_3103 = slice_3096 * slice_3102;
assign mul_3859 = slice_3856 * slice_3858;
assign addW_4615 = slice_4595 + slice_4577;
assign mul_708 = slice_706 * slice_707;
assign mul_5371 = slice_5369 * slice_5370;
assign addW_1464 = slice_1444 + slice_1402;
assign addW_6127 = slice_6122 + slice_6118;
assign slice_2220 = addW_2219[33:18];
assign mulnw_6883 = slice_6882 * slice_6879;
assign mul_2976 = slice_2970 * slice_2972;
assign mul_3732 = slice_3728 * slice_3731;
assign slice_4488 = slice_4487[63:32];
assign slice_581 = slice_580[32:16];
assign mulnw_5244 = slice_5242 * slice_5243;
assign slice_1337 = slice_1315[7:0];
assign addW_6000 = slice_5995 + slice_5990;
assign slice_2093 = slice_2092[31:18];
assign slice_6756 = slice_6735[16:8];
assign addW_2849 = slice_2844 + slice_2841;
assign mul_7512 = slice_7506 * slice_7508;
assign subW_3605 = subW_3604 - mul_3598;
assign add_4361 = lsl_4359 + mul_4360;
assign add_454 = lsl_452 + mul_453;
assign concat_5117 = {addW_5115,slice_5116};
assign add_1210 = lsl_1208 + mul_1209;
assign mul_5873 = slice_5871 * slice_5872;
assign addW_1966 = slice_1961 + slice_1958;
assign add_6629 = lsl_6620 + add_6628;
assign slice_2722 = concat_2676[31:0];
assign subW_7385 = concat_7384 - concat_7346;
assign subW_3478 = subW_3477 - mul_3471;
assign mulnw_4234 = slice_4227 * slice_4233;
assign concat_327 = {addW_325,slice_326};
assign add_4990 = lsl_4981 + add_4989;
assign addW_1083 = concat_1055 + addW_1082;
assign concat_5746 = {mul_5741,slice_5745};
assign mulnw_1839 = slice_1838 * slice_1835;
assign mul_6502 = slice_6500 * slice_6501;
assign slice_2595 = addW_2594[32:16];
assign mulnw_7258 = slice_7257 * slice_7254;
assign addW_3351 = slice_3346 + slice_3343;
assign lsl_4107 = mulnw_4106 << 16;
assign add_200 = lsl_191 + add_199;
assign add_4863 = lsl_4854 + add_4862;
assign concat_956 = {addW_954,slice_955};
assign mul_5619 = slice_5617 * slice_5618;
assign slice_1712 = slice_1707[15:8];
assign add_6375 = lsl_6373 + mul_6374;
assign slice_2468 = addW_2426[32:0];
assign addW_7131 = slice_7126 + slice_7122;
assign mulnw_3224 = slice_3223 * slice_3220;
assign addW_3980 = slice_3975 + slice_3972;
assign subW_4736 = subW_4735 - mul_4729;
assign addW_829 = concat_801 + addW_828;
assign slice_5492 = slice_5474[15:8];
assign concat_1585 = {mul_1580,slice_1584};
assign subW_6248 = subW_6247 - concat_6204;
assign slice_2341 = addW_2255[64:0];
assign subW_7004 = concat_7003 - concat_6943;
assign slice_3097 = slice_3092[15:8];
assign slice_3853 = mul_3822[15:0];
assign slice_4609 = mul_4600[17:0];
assign slice_702 = addW_701[32:16];
assign slice_5365 = slice_5364[31:18];
assign subW_1458 = subW_1457 - mul_1451;
assign mul_6121 = slice_6118 * slice_6120;
assign addW_2214 = concat_2208 + subW_2213;
assign add_6877 = lsl_6868 + add_6876;
assign slice_2970 = slice_2948[7:0];
assign slice_3726 = slice_3639[63:0];
assign subW_4482 = subW_4481 - concat_4371;
assign slice_575 = addW_574[128:64];
assign slice_5238 = slice_5234[15:0];
assign add_1331 = lsl_1329 + mul_1330;
assign mul_5994 = slice_5990 * slice_5993;
assign addW_2087 = concat_2081 + subW_2086;
assign add_6750 = mulnw_6747 + mulnw_6749;
assign slice_2843 = slice_2838[17:0];
assign slice_7506 = slice_7484[7:0];
assign slice_3599 = mul_3598[35:18];
assign mulnw_4355 = slice_4354 * slice_4351;
assign mulnw_448 = slice_447 * slice_444;
assign addW_5111 = slice_5106 + slice_5103;
assign mulnw_1204 = slice_1203 * slice_1200;
assign slice_5867 = addW_5866[33:18];
assign slice_1960 = addW_1955[17:0];
assign slice_6623 = slice_6613[7:0];
assign addW_2716 = concat_2688 + addW_2715;
assign mul_7379 = addW_7377 * addW_7378;
assign slice_3472 = mul_3471[35:18];
assign slice_4228 = slice_4207[16:8];
assign addW_321 = slice_316 + slice_313;
assign slice_4984 = slice_4974[7:0];
assign add_1077 = mulnw_1074 + mulnw_1076;
assign slice_5740 = slice_5739[31:18];
assign concat_1833 = {mul_1828,slice_1832};
assign slice_6496 = addW_6495[33:18];
assign addW_2589 = concat_2583 + subW_2588;
assign add_7252 = lsl_7243 + add_7251;
assign slice_3345 = addW_3340[17:0];
assign mul_4101 = slice_4095 * slice_4097;
assign slice_194 = slice_168[7:0];
assign slice_4857 = slice_4847[7:0];
assign slice_950 = mul_919[15:0];
assign slice_5613 = addW_5612[129:65];
assign slice_1706 = slice_1698[15:0];
assign mulnw_6369 = slice_6368 * slice_6365;
assign add_2462 = lsl_2460 + mul_2461;
assign mul_7125 = slice_7122 * slice_7124;
assign concat_3218 = {mul_3213,slice_3217};
assign slice_3974 = addW_3969[17:0];
assign addW_67 = concat_61 + subW_66;
assign slice_4730 = mul_4729[35:18];
assign add_823 = mulnw_820 + mulnw_822;
assign mulnw_5486 = slice_5479 * slice_5485;
assign slice_1579 = slice_1578[32:16];
assign add_6242 = lsl_6233 + add_6241;
assign addW_2335 = concat_2314 + subW_2334;
assign mul_6998 = addW_6996 * addW_6997;
assign slice_3091 = slice_3084[15:0];
assign lsl_3847 = add_3846 << 8;
assign addW_4603 = slice_4598 + slice_4594;
assign addW_696 = concat_690 + subW_695;
assign subW_5359 = mul_5358 - mul_5350;
assign slice_1452 = mul_1451[35:18];
assign slice_6115 = mul_6084[15:0];
assign concat_2208 = {mul_2203,slice_2207};
assign slice_6871 = slice_6861[7:0];
assign add_2964 = lsl_2962 + mul_2963;
assign concat_3720 = {addW_3718,slice_3719};
assign subW_4476 = concat_4475 - concat_4415;
assign concat_569 = {addW_567,slice_568};
assign slice_5232 = slice_5231[32:16];
assign mulnw_1325 = slice_1324 * slice_1321;
assign slice_5988 = slice_5900[63:0];
assign concat_2081 = {mul_2076,slice_2080};
assign mulnw_6744 = slice_6742 * slice_6743;
assign concat_2837 = {addW_2835,slice_2836};
assign add_7500 = lsl_7498 + mul_7499;
assign slice_3593 = addW_3552[31:0];
assign add_4349 = lsl_4340 + add_4348;
assign concat_442 = {mul_437,slice_441};
assign slice_5105 = slice_5100[17:0];
assign add_1198 = lsl_1189 + add_1197;
assign addW_5861 = concat_5833 + addW_5860;
assign concat_1954 = {concat_1912,slice_1953};
assign slice_6617 = slice_6607[16:8];
assign add_2710 = mulnw_2707 + mulnw_2709;
assign slice_7373 = addW_7369[17:0];
assign slice_3466 = slice_3465[63:32];
assign add_4222 = mulnw_4219 + mulnw_4221;
assign slice_315 = slice_308[17:0];
assign slice_4978 = slice_4969[16:8];
assign mulnw_1071 = slice_1069 * slice_1070;
assign addW_5734 = concat_5706 + addW_5733;
assign slice_1827 = addW_1826[32:16];
assign addW_6490 = concat_6484 + subW_6489;
assign concat_2583 = {mul_2578,slice_2582};
assign slice_7246 = slice_7236[7:0];
assign concat_3339 = {concat_3297,slice_3338};
assign slice_4095 = slice_4081[7:0];
assign slice_188 = slice_170[15:8];
assign slice_4851 = slice_4841[16:8];
assign lsl_944 = add_943 << 8;
assign concat_5607 = {concat_5341,slice_5606};
assign addW_1700 = slice_873 + slice_28;
assign add_6363 = lsl_6354 + add_6362;
assign mulnw_2456 = slice_2455 * slice_2452;
assign slice_7119 = mul_7110[17:0];
assign slice_3212 = addW_3211[32:16];
assign concat_3968 = {concat_3948,slice_3967};
assign concat_61 = {mul_56,slice_60};
assign addW_4724 = slice_4704 + slice_4664;
assign mulnw_817 = slice_815 * slice_816;
assign slice_5480 = slice_5475[15:8];
assign concat_1573 = {concat_1486,slice_1572};
assign slice_6236 = slice_6210[7:0];
assign subW_2329 = subW_2328 - mul_2322;
assign slice_6992 = addW_6988[17:0];
assign slice_3085 = slice_3084[32:16];
assign lsl_3841 = mulnw_3840 << 16;
assign mul_4597 = slice_4594 * slice_4596;
assign concat_690 = {mul_685,slice_689};
assign mul_5353 = slice_5351 * slice_5352;
assign slice_1446 = slice_1405[31:0];
assign lsl_6109 = add_6108 << 8;
assign slice_2202 = slice_2201[31:18];
assign slice_6865 = slice_6856[16:8];
assign mulnw_2958 = slice_2957 * slice_2954;
assign mul_3714 = slice_3708 * slice_3710;
assign mul_4470 = addW_4468 * addW_4469;
assign slice_563 = concat_539[31:0];
assign slice_5226 = concat_5180[31:0];
assign concat_1319 = {mul_1314,slice_1318};
assign concat_5982 = {addW_5980,slice_5981};
assign slice_2075 = slice_2074[31:18];
assign slice_6738 = slice_6734[15:0];
assign addW_2831 = slice_2826 + slice_2823;
assign mulnw_7494 = slice_7493 * slice_7490;
assign addW_3587 = add_3573 + add_3586;
assign slice_4343 = slice_4333[7:0];
assign slice_436 = addW_435[32:16];
assign concat_5099 = {addW_5097,slice_5098};
assign slice_1192 = slice_1182[7:0];
assign add_5855 = mulnw_5852 + mulnw_5854;
assign add_1948 = lsl_1939 + add_1947;
assign mul_6611 = slice_6607 * slice_6610;
assign mulnw_2704 = slice_2702 * slice_2703;
assign addW_7367 = slice_7347 + slice_7305;
assign slice_3460 = concat_3414[31:0];
assign mulnw_4216 = slice_4214 * slice_4215;
assign slice_309 = slice_308[31:18];
assign mul_4972 = slice_4969 * slice_4971;
assign lsl_1065 = add_1064 << 8;
assign add_5728 = mulnw_5725 + mulnw_5727;
assign concat_1821 = {addW_1819,slice_1820};
assign concat_6484 = {mul_6479,slice_6483};
assign slice_2577 = slice_2576[31:18];
assign slice_7240 = slice_7231[16:8];
assign add_3333 = lsl_3324 + add_3332;
assign slice_4089 = mul_4088[31:16];
assign mulnw_182 = slice_175 * slice_181;
assign mul_4845 = slice_4841 * slice_4844;
assign lsl_938 = mulnw_937 << 16;
assign subW_5601 = concat_5600 - concat_5428;
assign slice_6357 = slice_6347[7:0];
assign add_2450 = lsl_2441 + add_2449;
assign addW_7113 = slice_7108 + slice_7103;
assign concat_3206 = {addW_3204,slice_3205};
assign subW_3962 = mul_3961 - mul_3953;
assign slice_55 = slice_54[31:18];
assign slice_4718 = mul_4709[17:0];
assign lsl_811 = add_810 << 8;
assign slice_5474 = addW_5469[15:0];
assign subW_1567 = concat_1566 - concat_1506;
assign slice_6230 = slice_6212[15:8];
assign slice_2323 = mul_2322[35:18];
assign addW_6986 = slice_6944 + slice_6903;
assign concat_3079 = {addW_3077,slice_3078};
assign mul_3835 = slice_3829 * slice_3831;
assign slice_4591 = mul_4582[17:0];
assign slice_684 = slice_683[31:18];
assign slice_5347 = slice_5346[127:64];
assign addW_1440 = add_1426 + add_1439;
assign lsl_6103 = mulnw_6102 << 16;
assign addW_2196 = concat_2168 + addW_2195;
assign mul_6859 = slice_6856 * slice_6858;
assign concat_2952 = {mul_2947,slice_2951};
assign slice_3708 = slice_3686[7:0];
assign slice_4464 = addW_4460[17:0];
assign addW_557 = concat_551 + subW_556;
assign addW_5220 = concat_5192 + addW_5219;
assign slice_1313 = slice_1312[32:16];
assign mul_5976 = slice_5970 * slice_5972;
assign concat_2069 = {addW_2067,slice_2068};
assign slice_6732 = addW_6731[257:129];
assign slice_2825 = slice_2818[17:0];
assign concat_7488 = {mul_7483,slice_7487};
assign mulnw_3581 = slice_3574 * slice_3580;
assign slice_4337 = slice_4328[16:8];
assign concat_430 = {addW_428,slice_429};
assign mul_5093 = slice_5087 * slice_5089;
assign slice_1186 = slice_1177[16:8];
assign mulnw_5849 = slice_5847 * slice_5848;
assign slice_1942 = slice_1916[7:0];
assign addW_6605 = slice_6518 + slice_6432;
assign lsl_2698 = add_2697 << 8;
assign subW_7361 = subW_7360 - mul_7354;
assign addW_3454 = concat_3426 + addW_3453;
assign slice_4210 = slice_4206[15:0];
assign addW_303 = concat_211 + subW_302;
assign slice_4966 = mul_4935[15:0];
assign lsl_1059 = mulnw_1058 << 16;
assign mulnw_5722 = slice_5720 * slice_5721;
assign addW_1815 = slice_1810 + slice_1807;
assign slice_6478 = slice_6477[31:18];
assign addW_2571 = concat_2565 + subW_2570;
assign mul_7234 = slice_7231 * slice_7233;
assign slice_3327 = slice_3301[7:0];
assign slice_4083 = addW_4082[65:33];
assign slice_176 = slice_171[15:8];
assign slice_4839 = addW_4752[64:0];
assign mul_932 = slice_926 * slice_928;
assign concat_5595 = {addW_5593,slice_5594};
assign addW_1688 = concat_1399 + subW_1687;
assign slice_6351 = slice_6341[16:8];
assign slice_2444 = slice_2434[7:0];
assign mul_7107 = slice_7103 * slice_7106;
assign addW_3200 = slice_3195 + slice_3192;
assign mul_3956 = slice_3954 * slice_3955;
assign addW_49 = concat_41 + subW_48;
assign addW_4712 = slice_4707 + slice_4703;
assign lsl_805 = mulnw_804 << 16;
assign concat_5468 = {concat_5448,slice_5467};
assign add_1561 = lsl_1559 + mul_1560;
assign mulnw_6224 = slice_6217 * slice_6223;
assign addW_2317 = slice_2297 + slice_2257;
assign addW_6980 = add_6966 + add_6979;
assign slice_3073 = concat_3049[31:0];
assign slice_3829 = slice_3815[7:0];
assign addW_4585 = slice_4580 + slice_4575;
assign addW_678 = concat_672 + subW_677;
assign concat_5341 = {addW_5339,slice_5340};
assign mulnw_1434 = slice_1427 * slice_1433;
assign mul_6097 = slice_6091 * slice_6093;
assign add_2190 = mulnw_2187 + mulnw_2189;
assign slice_6853 = concat_6852[63:32];
assign slice_2946 = addW_2945[32:16];
assign add_3702 = lsl_3700 + mul_3701;
assign addW_4458 = slice_4416 + slice_4375;
assign concat_551 = {mul_546,slice_550};
assign add_5214 = mulnw_5211 + mulnw_5213;
assign concat_1307 = {concat_1220,slice_1306};
assign slice_5970 = slice_5948[7:0];
assign slice_2063 = mul_2032[15:0];
assign addW_6726 = slice_5899 + slice_5053;
assign slice_2819 = slice_2818[31:18];
assign slice_7482 = slice_7481[32:16];
assign slice_3575 = slice_3554[16:8];
assign mul_4331 = slice_4328 * slice_4330;
assign addW_424 = slice_419 + slice_416;
assign slice_5087 = slice_5065[7:0];
assign mul_1180 = slice_1177 * slice_1179;
assign lsl_5843 = add_5842 << 8;
assign slice_1936 = slice_1918[15:8];
assign subW_6599 = subW_6598 - concat_6555;
assign lsl_2692 = mulnw_2691 << 16;
assign slice_7355 = mul_7354[35:18];
assign add_3448 = mulnw_3445 + mulnw_3447;
assign slice_4204 = addW_4203[256:128];
assign subW_297 = subW_296 - concat_273;
assign lsl_4960 = add_4959 << 8;
assign mul_1053 = slice_1051 * slice_1052;
assign lsl_5716 = add_5715 << 8;
assign slice_1809 = slice_1804[17:0];
assign addW_6472 = concat_6444 + addW_6471;
assign concat_2565 = {mul_2560,slice_2564};
assign slice_7228 = mul_7197[15:0];
assign slice_3321 = slice_3303[15:8];
assign slice_4077 = concat_4076[127:64];
assign slice_170 = addW_165[15:0];
assign concat_4833 = {addW_4831,slice_4832};
assign slice_926 = slice_913[7:0];
assign addW_5589 = slice_5584 + slice_5581;
assign subW_1682 = subW_1681 - concat_1571;
assign mul_6345 = slice_6341 * slice_6344;
assign slice_2438 = slice_2428[16:8];
assign slice_7101 = slice_7014[63:0];
assign slice_3194 = slice_3189[17:0];
assign slice_3950 = slice_3949[31:18];
assign mul_4706 = slice_4703 * slice_4705;
assign mul_799 = slice_797 * slice_798;
assign subW_5462 = mul_5461 - mul_5453;
assign mulnw_1555 = slice_1554 * slice_1551;
assign slice_6218 = slice_6213[15:8];
assign slice_2311 = mul_2302[17:0];
assign mulnw_6974 = slice_6967 * slice_6973;
assign addW_3067 = concat_3061 + subW_3066;
assign slice_3823 = mul_3822[31:16];
assign mul_4579 = slice_4575 * slice_4578;
assign concat_672 = {mul_667,slice_671};
assign slice_5335 = concat_5311[32:0];
assign slice_1428 = slice_1407[16:8];
assign slice_6091 = slice_6077[7:0];
assign mulnw_2184 = slice_2182 * slice_2183;
assign mul_6847 = addW_6845 * addW_6846;
assign concat_2940 = {addW_2938,slice_2939};
assign concat_7603 = {addW_7601,slice_7602};
assign mulnw_3696 = slice_3695 * slice_3692;
assign addW_4452 = add_4438 + add_4451;
assign slice_545 = addW_544[33:18];
assign mulnw_5208 = slice_5206 * slice_5207;
assign subW_1301 = concat_1300 - concat_1240;
assign add_5964 = lsl_5962 + mul_5963;
assign lsl_2057 = add_2056 << 8;
assign slice_6720 = concat_6428[127:0];
assign addW_2813 = concat_2725 + subW_2812;
assign concat_7476 = {concat_7389,slice_7475};
assign add_3569 = mulnw_3566 + mulnw_3568;
assign slice_4325 = concat_4324[63:32];
assign slice_418 = slice_413[17:0];
assign add_5081 = lsl_5079 + mul_5080;
assign slice_1174 = concat_1173[63:32];
assign lsl_5837 = mulnw_5836 << 16;
assign mulnw_1930 = slice_1923 * slice_1929;
assign add_6593 = lsl_6584 + add_6592;
assign mul_2686 = slice_2684 * slice_2685;
assign slice_7349 = slice_7308[31:0];
assign mulnw_3442 = slice_3440 * slice_3441;
assign addW_4198 = slice_3373 + slice_2549;
assign subW_291 = mul_290 - mul_282;
assign lsl_4954 = mulnw_4953 << 16;
assign addW_1047 = slice_960 + slice_875;
assign lsl_5710 = mulnw_5709 << 16;
assign concat_1803 = {addW_1801,slice_1802};
assign add_6466 = mulnw_6463 + mulnw_6465;
assign slice_2559 = slice_2558[31:18];
assign lsl_7222 = add_7221 << 8;
assign mulnw_3315 = slice_3308 * slice_3314;
assign concat_4071 = {addW_4069,slice_4070};
assign concat_164 = {concat_144,slice_163};
assign addW_4827 = slice_4822 + slice_4819;
assign slice_920 = mul_919[31:16];
assign slice_5583 = addW_5578[17:0];
assign subW_1676 = concat_1675 - concat_1615;
assign addW_6339 = slice_6252 + slice_6166;
assign mul_2432 = slice_2428 * slice_2431;
assign concat_7095 = {addW_7093,slice_7094};
assign concat_3188 = {addW_3186,slice_3187};
assign add_3944 = lsl_3935 + add_3943;
assign slice_37 = slice_31[17:0];
assign slice_4700 = mul_4669[15:0];
assign slice_793 = slice_792[32:16];
assign mul_5456 = slice_5454 * slice_5455;
assign add_1549 = lsl_1540 + add_1548;
assign slice_6212 = addW_6207[15:0];
assign addW_2305 = slice_2300 + slice_2296;
assign slice_6968 = slice_6947[16:8];
assign concat_3061 = {mul_3056,slice_3060};
assign slice_3817 = addW_3816[64:32];
assign slice_4573 = slice_4486[63:0];
assign slice_666 = slice_665[31:18];
assign addW_5329 = concat_5323 + subW_5328;
assign add_1422 = mulnw_1419 + mulnw_1421;
assign slice_6085 = mul_6084[31:16];
assign lsl_2178 = add_2177 << 8;
assign slice_6841 = slice_6837[17:0];
assign addW_2934 = slice_2929 + slice_2926;
assign slice_7597 = concat_6721[255:0];
assign concat_3690 = {mul_3685,slice_3689};
assign mulnw_4446 = slice_4439 * slice_4445;
assign concat_539 = {addW_537,slice_538};
assign lsl_5202 = add_5201 << 8;
assign add_1295 = lsl_1293 + mul_1294;
assign mulnw_5958 = slice_5957 * slice_5954;
assign lsl_2051 = mulnw_2050 << 16;
assign addW_6714 = concat_6604 + subW_6713;
assign subW_2807 = subW_2806 - concat_2785;
assign subW_7470 = concat_7469 - concat_7431;
assign mulnw_3563 = slice_3561 * slice_3562;
assign mul_4319 = addW_4317 * addW_4318;
assign concat_412 = {addW_410,slice_411};
assign mulnw_5075 = slice_5074 * slice_5071;
assign mul_1168 = addW_1166 * addW_1167;
assign mul_5831 = slice_5829 * slice_5830;
assign slice_1924 = slice_1919[15:8];
assign slice_6587 = slice_6561[7:0];
assign slice_2680 = addW_2679[32:16];
assign addW_7343 = add_7329 + add_7342;
assign lsl_3436 = add_3435 << 8;
assign subW_4192 = subW_4191 - concat_3902;
assign mul_285 = slice_283 * slice_284;
assign mul_4948 = slice_4942 * slice_4944;
assign concat_1041 = {addW_1039,slice_1040};
assign mul_5704 = slice_5702 * slice_5703;
assign addW_1797 = slice_1792 + slice_1789;
assign mulnw_6460 = slice_6458 * slice_6459;
assign slice_2553 = slice_2552[31:18];
assign lsl_7216 = mulnw_7215 << 16;
assign slice_3309 = slice_3304[15:8];
assign mul_4065 = slice_4059 * slice_4061;
assign subW_158 = mul_157 - mul_149;
assign slice_4821 = addW_4816[17:0];
assign addW_914 = slice_894 + slice_876;
assign concat_5577 = {concat_5557,slice_5576};
assign mul_1670 = addW_1668 * addW_1669;
assign subW_6333 = subW_6332 - concat_6289;
assign addW_2426 = slice_2338 + slice_2252;
assign addW_7089 = slice_7084 + slice_7081;
assign addW_3182 = slice_3177 + slice_3174;
assign slice_3938 = slice_3912[7:0];
assign slice_31 = slice_30[63:32];
assign lsl_4694 = add_4693 << 8;
assign add_787 = lsl_778 + add_786;
assign slice_5450 = slice_5449[31:18];
assign slice_1543 = slice_1533[7:0];
assign concat_6206 = {concat_6186,slice_6205};
assign mul_2299 = slice_2296 * slice_2298;
assign add_6962 = mulnw_6959 + mulnw_6961;
assign slice_3055 = addW_3054[33:18];
assign slice_3811 = concat_3810[127:64];
assign concat_4567 = {addW_4565,slice_4566};
assign concat_660 = {addW_658,slice_659};
assign concat_5323 = {mul_5318,slice_5322};
assign mulnw_1416 = slice_1414 * slice_1415;
assign slice_6079 = addW_6078[64:32];
assign lsl_2172 = mulnw_2171 << 16;
assign slice_6835 = slice_6815[31:0];
assign slice_2928 = slice_2923[17:0];
assign addW_7591 = concat_7301 + subW_7590;
assign slice_3684 = addW_3683[32:16];
assign slice_4440 = slice_4419[16:8];
assign addW_533 = slice_528 + slice_525;
assign lsl_5196 = mulnw_5195 << 16;
assign mulnw_1289 = slice_1288 * slice_1285;
assign concat_5952 = {mul_5947,slice_5951};
assign mul_2045 = slice_2039 * slice_2041;
assign subW_6708 = subW_6707 - concat_6686;
assign subW_2801 = mul_2800 - mul_2792;
assign mul_7464 = addW_7462 * addW_7463;
assign slice_3557 = slice_3553[15:0];
assign slice_4313 = slice_4309[17:0];
assign addW_406 = slice_401 + slice_398;
assign concat_5069 = {mul_5064,slice_5068};
assign slice_1162 = slice_1158[17:0];
assign slice_5825 = slice_5824[32:16];
assign slice_1918 = slice_1913[15:0];
assign slice_6581 = slice_6563[15:8];
assign addW_2674 = concat_2668 + subW_2673;
assign mulnw_7337 = slice_7330 * slice_7336;
assign lsl_3430 = mulnw_3429 << 16;
assign subW_4186 = concat_4185 - concat_3991;
assign slice_279 = addW_278[33:18];
assign slice_4942 = slice_4928[7:0];
assign slice_1035 = mul_1004[15:0];
assign slice_5698 = addW_5612[64:0];
assign slice_1791 = slice_1785[17:0];
assign lsl_6454 = add_6453 << 8;
assign concat_2547 = {addW_2545,slice_2546};
assign mul_7210 = slice_7204 * slice_7206;
assign slice_3303 = slice_3298[15:0];
assign slice_4059 = slice_4037[7:0];
assign mul_152 = slice_150 * slice_151;
assign concat_4815 = {concat_4795,slice_4814};
assign slice_908 = mul_899[17:0];
assign subW_5571 = mul_5570 - mul_5562;
assign slice_1664 = addW_1660[17:0];
assign add_6327 = lsl_6318 + add_6326;
assign addW_2420 = concat_2399 + subW_2419;
assign slice_7083 = addW_7078[17:0];
assign slice_3176 = slice_3170[17:0];
assign slice_3932 = slice_3914[15:8];
assign slice_25 = slice_22[31:18];
assign lsl_4688 = mulnw_4687 << 16;
assign slice_781 = slice_755[7:0];
assign subW_5444 = mul_5443 - mul_5435;
assign slice_1537 = slice_1528[16:8];
assign subW_6200 = mul_6199 - mul_6191;
assign slice_2293 = mul_2262[15:0];
assign mulnw_6956 = slice_6954 * slice_6955;
assign concat_3049 = {addW_3047,slice_3048};
assign concat_3805 = {addW_3803,slice_3804};
assign mul_4561 = slice_4555 * slice_4557;
assign slice_654 = mul_645[17:0];
assign slice_5317 = addW_5316[33:18];
assign slice_1410 = slice_1406[15:0];
assign slice_6073 = concat_6072[127:64];
assign mul_2166 = slice_2164 * slice_2165;
assign mul_6829 = addW_6827 * addW_6828;
assign concat_2922 = {addW_2920,slice_2921};
assign subW_7585 = subW_7584 - concat_7474;
assign concat_3678 = {addW_3676,slice_3677};
assign add_4434 = mulnw_4431 + mulnw_4433;
assign slice_527 = slice_522[17:0];
assign mul_5190 = slice_5188 * slice_5189;
assign add_1283 = lsl_1274 + add_1282;
assign slice_5946 = addW_5945[32:16];
assign slice_2039 = slice_2026[7:0];
assign subW_6702 = mul_6701 - mul_6693;
assign mul_2795 = slice_2793 * slice_2794;
assign slice_7458 = addW_7454[17:0];
assign slice_3551 = slice_3550[32:16];
assign slice_4307 = slice_4287[31:0];
assign slice_400 = slice_394[17:0];
assign slice_5063 = slice_5062[32:16];
assign slice_1156 = slice_1135[31:0];
assign add_5819 = lsl_5810 + add_5818;
assign concat_1912 = {addW_1910,slice_1911};
assign mulnw_6575 = slice_6568 * slice_6574;
assign concat_2668 = {mul_2663,slice_2667};
assign slice_7331 = slice_7310[16:8];
assign mul_3424 = slice_3422 * slice_3423;
assign concat_4180 = {addW_4178,slice_4179};
assign concat_273 = {addW_271,slice_272};
assign slice_4936 = mul_4935[31:16];
assign lsl_1029 = add_1028 << 8;
assign addW_5692 = concat_5671 + subW_5691;
assign slice_1785 = slice_1784[63:32];
assign lsl_6448 = mulnw_6447 << 16;
assign slice_2541 = concat_2246[127:0];
assign slice_7204 = slice_7190[7:0];
assign concat_3297 = {addW_3295,slice_3296};
assign add_4053 = lsl_4051 + mul_4052;
assign slice_146 = slice_145[31:18];
assign subW_4809 = mul_4808 - mul_4800;
assign addW_902 = slice_897 + slice_893;
assign mul_5565 = slice_5563 * slice_5564;
assign addW_1658 = slice_1616 + slice_1575;
assign slice_6321 = slice_6295[7:0];
assign subW_2414 = subW_2413 - mul_2407;
assign concat_7077 = {concat_7057,slice_7076};
assign slice_3170 = slice_3169[63:32];
assign mulnw_3926 = slice_3919 * slice_3925;
assign slice_19 = slice_16[127:64];
assign mul_4682 = slice_4676 * slice_4678;
assign slice_775 = slice_757[15:8];
assign mul_5438 = slice_5436 * slice_5437;
assign mul_1531 = slice_1528 * slice_1530;
assign mul_6194 = slice_6192 * slice_6193;
assign lsl_2287 = add_2286 << 8;
assign slice_6950 = slice_6946[15:0];
assign addW_3043 = slice_3038 + slice_3035;
assign mul_3799 = slice_3793 * slice_3795;
assign slice_4555 = slice_4533[7:0];
assign addW_648 = slice_643 + slice_639;
assign concat_5311 = {addW_5309,slice_5310};
assign addW_1404 = slice_1138 + slice_874;
assign concat_6067 = {addW_6065,slice_6066};
assign addW_2160 = slice_2073 + slice_1988;
assign slice_6823 = slice_6819[17:0];
assign addW_2916 = slice_2911 + slice_2908;
assign subW_7579 = concat_7578 - concat_7518;
assign addW_3672 = slice_3667 + slice_3664;
assign mulnw_4428 = slice_4426 * slice_4427;
assign concat_521 = {addW_519,slice_520};
assign slice_5184 = addW_5183[32:16];
assign slice_1277 = slice_1267[7:0];
assign concat_5940 = {addW_5938,slice_5939};
assign slice_2033 = mul_2032[31:16];
assign mul_6696 = slice_6694 * slice_6695;
assign slice_2789 = addW_2788[33:18];
assign addW_7452 = slice_7432 + slice_7391;
assign slice_3545 = concat_3499[31:0];
assign mul_4301 = addW_4299 * addW_4300;
assign slice_394 = slice_393[63:32];
assign slice_5057 = slice_5056[32:16];
assign mul_1150 = addW_1148 * addW_1149;
assign slice_5813 = slice_5787[7:0];
assign mul_1906 = slice_1900 * slice_1902;
assign slice_6569 = slice_6564[15:8];
assign slice_2662 = slice_2661[31:18];
assign add_7325 = mulnw_7322 + mulnw_7324;
assign slice_3418 = addW_3417[32:16];
assign addW_4174 = slice_4169 + slice_4166;
assign addW_267 = slice_262 + slice_259;
assign slice_4930 = addW_4929[65:33];
assign lsl_1023 = mulnw_1022 << 16;
assign subW_5686 = subW_5685 - mul_5679;
assign subW_1779 = concat_1778 - concat_1740;
assign mul_6442 = slice_6440 * slice_6441;
assign addW_2535 = concat_2424 + subW_2534;
assign slice_7198 = mul_7197[31:16];
assign mul_3291 = slice_3285 * slice_3287;
assign mulnw_4047 = slice_4046 * slice_4043;
assign subW_140 = mul_139 - mul_131;
assign mul_4803 = slice_4801 * slice_4802;
assign mul_896 = slice_893 * slice_895;
assign slice_5559 = slice_5558[31:18];
assign addW_1652 = add_1638 + add_1651;
assign slice_6315 = slice_6297[15:8];
assign slice_2408 = mul_2407[35:18];
assign subW_7071 = mul_7070 - mul_7062;
assign subW_3164 = concat_3163 - concat_3125;
assign slice_3920 = slice_3915[15:8];
assign slice_13 = slice_10[511:256];
assign slice_4676 = slice_4662[7:0];
assign mulnw_769 = slice_762 * slice_768;
assign slice_5432 = slice_5346[63:0];
assign slice_1525 = concat_1524[63:32];
assign slice_6188 = slice_6187[31:18];
assign lsl_2281 = mulnw_2280 << 16;
assign slice_6944 = addW_6902[32:0];
assign slice_3037 = slice_3032[17:0];
assign slice_3793 = slice_3771[7:0];
assign add_4549 = lsl_4547 + mul_4548;
assign mul_642 = slice_639 * slice_641;
assign mul_5305 = slice_5299 * slice_5301;
assign slice_1398 = concat_1397[255:128];
assign mul_6061 = slice_6055 * slice_6057;
assign concat_2154 = {addW_2152,slice_2153};
assign slice_6817 = slice_6816[31:18];
assign slice_2910 = slice_2904[17:0];
assign mul_7573 = addW_7571 * addW_7572;
assign slice_3666 = slice_3661[17:0];
assign slice_4422 = slice_4418[15:0];
assign mul_515 = slice_509 * slice_511;
assign addW_5178 = concat_5172 + subW_5177;
assign slice_1271 = slice_1262[16:8];
assign addW_5934 = slice_5929 + slice_5926;
assign addW_2027 = slice_2007 + slice_1989;
assign slice_6690 = addW_6689[33:18];
assign addW_2783 = concat_2777 + subW_2782;
assign subW_7446 = subW_7445 - mul_7439;
assign addW_3539 = concat_3511 + addW_3538;
assign slice_4295 = slice_4291[17:0];
assign subW_388 = concat_387 - concat_327;
assign slice_1144 = slice_1140[17:0];
assign slice_5807 = slice_5789[15:8];
assign slice_1900 = slice_1878[7:0];
assign slice_6563 = addW_6558[15:0];
assign addW_2656 = concat_2650 + subW_2655;
assign mulnw_7319 = slice_7317 * slice_7318;
assign addW_3412 = concat_3406 + subW_3411;
assign slice_4168 = addW_4163[17:0];
assign slice_261 = slice_256[17:0];
assign slice_4924 = concat_4923[129:65];
assign mul_1017 = slice_1011 * slice_1013;
assign slice_5680 = mul_5679[35:18];
assign mul_1773 = addW_1771 * addW_1772;
assign slice_6436 = addW_6435[128:64];
assign subW_2529 = subW_2528 - concat_2507;
assign slice_7192 = addW_7191[65:33];
assign slice_3285 = slice_3263[7:0];
assign concat_4041 = {mul_4036,slice_4040};
assign mul_134 = slice_132 * slice_133;
assign slice_4797 = slice_4796[31:18];
assign slice_890 = mul_881[17:0];
assign add_5553 = lsl_5544 + add_5552;
assign mulnw_1646 = slice_1639 * slice_1645;
assign mulnw_6309 = slice_6302 * slice_6308;
assign addW_2402 = slice_2382 + slice_2342;
assign mul_7065 = slice_7063 * slice_7064;
assign mul_3158 = addW_3156 * addW_3157;
assign slice_3914 = slice_3907[15:0];
assign slice_4670 = mul_4669[31:16];
assign slice_763 = slice_758[15:8];
assign addW_5426 = concat_5383 + subW_5425;
assign mul_1519 = addW_1517 * addW_1518;
assign subW_6182 = mul_6181 - mul_6173;
assign mul_2275 = slice_2269 * slice_2271;
assign add_6938 = lsl_6936 + mul_6937;
assign concat_3031 = {addW_3029,slice_3030};
assign add_3787 = lsl_3785 + mul_3786;
assign mulnw_4543 = slice_4542 * slice_4539;
assign slice_636 = concat_635[63:32];
assign slice_5299 = slice_5277[7:0];
assign concat_1392 = {addW_1390,slice_1391};
assign slice_6055 = slice_6033[7:0];
assign slice_2148 = mul_2117[15:0];
assign subW_6811 = subW_6810 - concat_6789;
assign slice_2904 = slice_2903[63:32];
assign slice_7567 = addW_7563[17:0];
assign concat_3660 = {addW_3658,slice_3659};
assign slice_4416 = addW_4374[32:0];
assign slice_509 = slice_487[7:0];
assign concat_5172 = {mul_5167,slice_5171};
assign mul_1265 = slice_1262 * slice_1264;
assign slice_5928 = slice_5923[17:0];
assign slice_2021 = mul_2012[17:0];
assign addW_6684 = concat_6656 + addW_6683;
assign concat_2777 = {mul_2772,slice_2776};
assign slice_7440 = mul_7439[35:18];
assign add_3533 = mulnw_3530 + mulnw_3532;
assign slice_4289 = slice_4288[31:18];
assign add_382 = lsl_380 + mul_381;
assign addW_5045 = concat_4197 + subW_5044;
assign slice_1138 = slice_873[127:0];
assign mulnw_5801 = slice_5794 * slice_5800;
assign add_1894 = lsl_1892 + mul_1893;
assign concat_6557 = {concat_6537,slice_6556};
assign concat_2650 = {mul_2645,slice_2649};
assign slice_7313 = slice_7309[15:0];
assign concat_3406 = {mul_3401,slice_3405};
assign concat_4162 = {concat_4120,slice_4161};
assign concat_255 = {addW_253,slice_254};
assign concat_4918 = {addW_4916,slice_4917};
assign slice_1011 = slice_998[7:0];
assign addW_5674 = slice_5654 + slice_5614;
assign slice_1767 = addW_1763[17:0];
assign concat_6430 = {concat_6164,slice_6429};
assign subW_2523 = mul_2522 - mul_2514;
assign slice_7186 = concat_7185[127:64];
assign add_3279 = lsl_3277 + mul_3278;
assign slice_4035 = addW_4034[32:16];
assign slice_128 = slice_29[63:0];
assign add_4791 = lsl_4782 + add_4790;
assign addW_884 = slice_879 + slice_872;
assign slice_5547 = slice_5521[7:0];
assign slice_1640 = slice_1619[16:8];
assign slice_6303 = slice_6298[15:8];
assign slice_2396 = mul_2387[17:0];
assign slice_7059 = slice_7058[31:18];
assign slice_3152 = addW_3148[17:0];
assign slice_3908 = slice_3907[32:16];
assign slice_4664 = addW_4663[64:32];
assign slice_757 = slice_751[15:0];
assign addW_5420 = add_5406 + add_5419;
assign slice_1513 = slice_1509[17:0];
assign mul_6176 = slice_6174 * slice_6175;
assign slice_2269 = slice_2254[7:0];
assign mulnw_6932 = slice_6931 * slice_6928;
assign mul_3025 = slice_3019 * slice_3021;
assign mulnw_3781 = slice_3780 * slice_3777;
assign concat_4537 = {mul_4532,slice_4536};
assign mul_630 = addW_628 * addW_629;
assign add_5293 = lsl_5291 + mul_5292;
assign slice_1386 = mul_1377[17:0];
assign add_6049 = lsl_6047 + mul_6048;
assign lsl_2142 = add_2141 << 8;
assign subW_6805 = mul_6804 - mul_6796;
assign subW_2898 = concat_2897 - concat_2837;
assign addW_7561 = slice_7519 + slice_7478;
assign addW_3654 = slice_3649 + slice_3646;
assign add_4410 = lsl_4408 + mul_4409;
assign add_503 = lsl_501 + mul_502;
assign slice_5166 = slice_5165[31:18];
assign slice_1259 = concat_1258[63:32];
assign concat_5922 = {addW_5920,slice_5921};
assign addW_2015 = slice_2010 + slice_2006;
assign add_6678 = mulnw_6675 + mulnw_6677;
assign slice_2771 = slice_2770[31:18];
assign slice_7434 = slice_7393[31:0];
assign mulnw_3527 = slice_3525 * slice_3526;
assign subW_4283 = subW_4282 - concat_4261;
assign mulnw_376 = slice_375 * slice_372;
assign subW_5039 = subW_5038 - concat_4749;
assign slice_1132 = concat_1041[63:0];
assign slice_5795 = slice_5790[15:8];
assign mulnw_1888 = slice_1887 * slice_1884;
assign subW_6551 = mul_6550 - mul_6542;
assign slice_2644 = slice_2643[31:18];
assign addW_7307 = slice_7018 + slice_6732;
assign slice_3400 = slice_3399[31:18];
assign add_4156 = lsl_4147 + add_4155;
assign mul_249 = slice_243 * slice_245;
assign addW_4912 = slice_4907 + slice_4904;
assign slice_1005 = mul_1004[31:16];
assign slice_5668 = mul_5659[17:0];
assign addW_1761 = slice_1741 + slice_1698;
assign subW_6424 = concat_6423 - concat_6251;
assign mul_2517 = slice_2515 * slice_2516;
assign concat_7180 = {addW_7178,slice_7179};
assign mulnw_3273 = slice_3272 * slice_3269;
assign concat_4029 = {addW_4027,slice_4028};
assign addW_122 = concat_71 + subW_121;
assign slice_4785 = slice_4759[7:0];
assign mul_878 = slice_872 * slice_877;
assign slice_5541 = slice_5523[15:8];
assign add_1634 = mulnw_1631 + mulnw_1633;
assign slice_6297 = addW_6292[15:0];
assign addW_2390 = slice_2385 + slice_2381;
assign add_7053 = lsl_7044 + add_7052;
assign addW_3146 = slice_3126 + slice_3084;
assign concat_3902 = {addW_3900,slice_3901};
assign slice_4658 = concat_4657[127:64];
assign slice_751 = addW_750[65:33];
assign mulnw_5414 = slice_5407 * slice_5413;
assign slice_1507 = slice_1487[31:0];
assign slice_6170 = slice_6169[127:64];
assign slice_2263 = mul_2262[31:16];
assign add_6926 = lsl_6917 + add_6925;
assign slice_3019 = slice_2997[7:0];
assign concat_3775 = {mul_3770,slice_3774};
assign slice_4531 = addW_4530[32:16];
assign slice_624 = slice_620[17:0];
assign mulnw_5287 = slice_5286 * slice_5283;
assign addW_1380 = slice_1375 + slice_1371;
assign mulnw_6043 = slice_6042 * slice_6039;
assign lsl_2136 = mulnw_2135 << 16;
assign mul_6799 = slice_6797 * slice_6798;
assign add_2892 = lsl_2890 + mul_2891;
assign addW_7555 = add_7541 + add_7554;
assign slice_3648 = slice_3641[17:0];
assign mulnw_4404 = slice_4403 * slice_4400;
assign mulnw_497 = slice_496 * slice_493;
assign addW_5160 = concat_5154 + subW_5159;
assign mul_1253 = addW_1251 * addW_1252;
assign addW_5916 = slice_5911 + slice_5908;
assign mul_2009 = slice_2006 * slice_2008;
assign mulnw_6672 = slice_6670 * slice_6671;
assign addW_2765 = concat_2737 + addW_2764;
assign addW_7428 = add_7414 + add_7427;
assign lsl_3521 = add_3520 << 8;
assign subW_4277 = mul_4276 - mul_4268;
assign add_370 = lsl_361 + add_369;
assign subW_5033 = concat_5032 - concat_4838;
assign addW_1126 = concat_1105 + subW_1125;
assign slice_5789 = slice_5783[15:0];
assign concat_1882 = {mul_1877,slice_1881};
assign mul_6545 = slice_6543 * slice_6544;
assign concat_2638 = {addW_2636,slice_2637};
assign concat_7301 = {concat_7013,slice_7300};
assign addW_3394 = concat_3388 + subW_3393;
assign slice_4150 = slice_4124[7:0];
assign slice_243 = slice_221[7:0];
assign slice_4906 = addW_4901[17:0];
assign addW_999 = slice_979 + slice_961;
assign addW_5662 = slice_5657 + slice_5653;
assign subW_1755 = subW_1754 - mul_1748;
assign concat_6418 = {addW_6416,slice_6417};
assign slice_2511 = addW_2510[33:18];
assign mul_7174 = slice_7168 * slice_7170;
assign concat_3267 = {mul_3262,slice_3266};
assign addW_4023 = slice_4018 + slice_4015;
assign addW_116 = add_102 + add_115;
assign slice_4779 = slice_4761[15:8];
assign slice_872 = slice_871[31:18];
assign mulnw_5535 = slice_5528 * slice_5534;
assign mulnw_1628 = slice_1626 * slice_1627;
assign concat_6291 = {concat_6271,slice_6290};
assign mul_2384 = slice_2381 * slice_2383;
assign slice_7047 = slice_7021[7:0];
assign subW_3140 = subW_3139 - mul_3133;
assign slice_3896 = concat_3872[31:0];
assign concat_4652 = {addW_4650,slice_4651};
assign concat_745 = {addW_743,slice_744};
assign slice_5408 = slice_5387[16:8];
assign mul_1501 = addW_1499 * addW_1500;
assign concat_6164 = {addW_6162,slice_6163};
assign slice_2257 = slice_2256[64:32];
assign slice_6920 = slice_6910[7:0];
assign add_3013 = lsl_3011 + mul_3012;
assign slice_3769 = addW_3768[32:16];
assign concat_4525 = {addW_4523,slice_4524};
assign slice_618 = slice_575[31:0];
assign concat_5281 = {mul_5276,slice_5280};
assign mul_1374 = slice_1371 * slice_1373;
assign concat_6037 = {mul_6032,slice_6036};
assign mul_2130 = slice_2124 * slice_2126;
assign slice_6793 = addW_6792[33:18];
assign mulnw_2886 = slice_2885 * slice_2882;
assign mulnw_7549 = slice_7542 * slice_7548;
assign slice_3642 = slice_3641[31:18];
assign add_4398 = lsl_4389 + add_4397;
assign concat_491 = {mul_486,slice_490};
assign concat_5154 = {mul_5149,slice_5153};
assign slice_1247 = slice_1243[17:0];
assign slice_5910 = slice_5902[17:0];
assign slice_2003 = mul_1994[17:0];
assign lsl_6666 = add_6665 << 8;
assign add_2759 = mulnw_2756 + mulnw_2758;
assign mulnw_7422 = slice_7415 * slice_7421;
assign lsl_3515 = mulnw_3514 << 16;
assign mul_4271 = slice_4269 * slice_4270;
assign slice_364 = slice_354[7:0];
assign concat_5027 = {addW_5025,slice_5026};
assign subW_1120 = subW_1119 - mul_1113;
assign slice_5783 = addW_5782[65:33];
assign slice_1876 = slice_1875[32:16];
assign slice_6539 = slice_6538[31:18];
assign slice_2632 = mul_2601[15:0];
assign subW_7295 = concat_7294 - concat_7100;
assign concat_3388 = {mul_3383,slice_3387};
assign slice_4144 = slice_4126[15:8];
assign add_237 = lsl_235 + mul_236;
assign concat_4900 = {concat_4880,slice_4899};
assign slice_993 = mul_984[17:0];
assign mul_5656 = slice_5653 * slice_5655;
assign slice_1749 = mul_1748[35:18];
assign addW_6412 = slice_6407 + slice_6404;
assign addW_2505 = concat_2477 + addW_2504;
assign slice_7168 = slice_7146[7:0];
assign slice_3261 = slice_3260[32:16];
assign slice_4017 = slice_4012[17:0];
assign mulnw_110 = slice_103 * slice_109;
assign mulnw_4773 = slice_4766 * slice_4772;
assign slice_866 = concat_569[127:0];
assign slice_5529 = slice_5524[15:8];
assign slice_1622 = slice_1618[15:0];
assign subW_6285 = mul_6284 - mul_6276;
assign slice_2378 = mul_2347[15:0];
assign slice_7041 = slice_7023[15:8];
assign slice_3134 = mul_3133[35:18];
assign addW_3890 = concat_3884 + subW_3889;
assign mul_4646 = slice_4640 * slice_4642;
assign slice_739 = mul_708[15:0];
assign add_5402 = mulnw_5399 + mulnw_5401;
assign slice_1495 = slice_1491[17:0];
assign slice_6158 = concat_6134[31:0];
assign addW_2251 = slice_1983 + slice_1696;
assign slice_6914 = slice_6904[16:8];
assign mulnw_3007 = slice_3006 * slice_3003;
assign concat_3763 = {addW_3761,slice_3762};
assign addW_4519 = slice_4514 + slice_4511;
assign add_612 = lsl_610 + mul_611;
assign slice_5275 = slice_5274[32:16];
assign slice_1368 = concat_1367[63:32];
assign slice_6031 = addW_6030[32:16];
assign slice_2124 = slice_2111[7:0];
assign addW_6787 = concat_6781 + subW_6786;
assign add_2880 = lsl_2871 + add_2879;
assign slice_7543 = slice_7522[16:8];
assign addW_3636 = concat_3548 + subW_3635;
assign slice_4392 = slice_4382[7:0];
assign slice_485 = slice_484[32:16];
assign slice_5148 = slice_5147[31:18];
assign slice_1241 = slice_1221[31:0];
assign slice_5904 = addW_5058[255:0];
assign addW_1997 = slice_1992 + slice_1986;
assign lsl_6660 = mulnw_6659 << 16;
assign mulnw_2753 = slice_2751 * slice_2752;
assign slice_7416 = slice_7395[16:8];
assign mul_3509 = slice_3507 * slice_3508;
assign slice_4265 = addW_4264[33:18];
assign slice_358 = slice_349[16:8];
assign addW_5021 = slice_5016 + slice_5013;
assign slice_1114 = mul_1113[35:18];
assign addW_5777 = concat_5756 + subW_5776;
assign concat_1870 = {concat_1783,slice_1869};
assign subW_6533 = mul_6532 - mul_6524;
assign lsl_2626 = add_2625 << 8;
assign concat_7289 = {addW_7287,slice_7288};
assign slice_3382 = slice_3381[31:18];
assign mulnw_4138 = slice_4131 * slice_4137;
assign mulnw_231 = slice_230 * slice_227;
assign subW_4894 = mul_4893 - mul_4885;
assign addW_987 = slice_982 + slice_978;
assign slice_5650 = mul_5619[15:0];
assign slice_1743 = slice_1702[31:0];
assign slice_6406 = addW_6401[17:0];
assign add_2499 = mulnw_2496 + mulnw_2498;
assign add_7162 = lsl_7160 + mul_7161;
assign concat_3255 = {concat_3168,slice_3254};
assign concat_4011 = {addW_4009,slice_4010};
assign slice_104 = slice_79[16:8];
assign slice_4767 = slice_4762[15:8];
assign addW_860 = concat_747 + subW_859;
assign slice_5523 = slice_5517[15:0];
assign slice_1616 = addW_1574[32:0];
assign mul_6279 = slice_6277 * slice_6278;
assign lsl_2372 = add_2371 << 8;
assign mulnw_7035 = slice_7028 * slice_7034;
assign slice_3128 = slice_3087[31:0];
assign concat_3884 = {mul_3879,slice_3883};
assign slice_4640 = slice_4618[7:0];
assign lsl_733 = add_732 << 8;
assign mulnw_5396 = slice_5394 * slice_5395;
assign slice_1489 = slice_1488[31:18];
assign addW_6152 = concat_6146 + subW_6151;
assign slice_2245 = concat_2154[63:0];
assign mul_6908 = slice_6904 * slice_6907;
assign concat_3001 = {mul_2996,slice_3000};
assign addW_3757 = slice_3752 + slice_3749;
assign slice_4513 = slice_4508[17:0];
assign mulnw_606 = slice_605 * slice_602;
assign addW_5269 = concat_5241 + addW_5268;
assign mul_1362 = addW_1360 * addW_1361;
assign concat_6025 = {addW_6023,slice_6024};
assign slice_2118 = mul_2117[31:16];
assign concat_6781 = {mul_6776,slice_6780};
assign slice_2874 = slice_2864[7:0];
assign add_7537 = mulnw_7534 + mulnw_7536;
assign subW_3630 = subW_3629 - concat_3608;
assign slice_4386 = slice_4376[16:8];
assign concat_479 = {concat_392,slice_478};
assign concat_5142 = {addW_5140,slice_5141};
assign mul_1235 = addW_1233 * addW_1234;
assign concat_5898 = {addW_5896,slice_5897};
assign mul_1991 = slice_1986 * slice_1990;
assign mul_6654 = slice_6652 * slice_6653;
assign lsl_2747 = add_2746 << 8;
assign add_7410 = mulnw_7407 + mulnw_7409;
assign slice_3503 = addW_3502[32:16];
assign addW_4259 = concat_4253 + subW_4258;
assign mul_352 = slice_349 * slice_351;
assign slice_5015 = addW_5010[17:0];
assign addW_1108 = slice_1088 + slice_1048;
assign subW_5771 = subW_5770 - mul_5764;
assign subW_1864 = concat_1863 - concat_1803;
assign mul_6527 = slice_6525 * slice_6526;
assign lsl_2620 = mulnw_2619 << 16;
assign addW_7283 = slice_7278 + slice_7275;
assign slice_3376 = slice_3375[63:32];
assign slice_4132 = slice_4127[15:8];
assign concat_225 = {mul_220,slice_224};
assign mul_4888 = slice_4886 * slice_4887;
assign mul_981 = slice_978 * slice_980;
assign lsl_5644 = add_5643 << 8;
assign addW_1737 = add_1723 + add_1736;
assign concat_6400 = {concat_6380,slice_6399};
assign mulnw_2493 = slice_2491 * slice_2492;
assign mulnw_7156 = slice_7155 * slice_7152;
assign subW_3249 = concat_3248 - concat_3188;
assign addW_4005 = slice_4000 + slice_3997;
assign add_98 = mulnw_95 + mulnw_97;
assign slice_4761 = slice_4754[15:0];
assign subW_854 = subW_853 - concat_831;
assign slice_5517 = addW_5516[64:32];
assign add_1610 = lsl_1608 + mul_1609;
assign slice_6273 = slice_6272[31:18];
assign lsl_2366 = mulnw_2365 << 16;
assign slice_7029 = slice_7024[15:8];
assign addW_3122 = add_3108 + add_3121;
assign slice_3878 = addW_3877[33:18];
assign add_4634 = lsl_4632 + mul_4633;
assign lsl_727 = mulnw_726 << 16;
assign slice_5390 = addW_5386[15:0];
assign subW_1483 = subW_1482 - concat_1461;
assign concat_6146 = {mul_6141,slice_6145};
assign addW_2239 = concat_2218 + subW_2238;
assign addW_6902 = slice_6815 + slice_6728;
assign slice_2995 = slice_2994[32:16];
assign slice_3751 = slice_3746[17:0];
assign concat_4507 = {addW_4505,slice_4506};
assign add_600 = lsl_591 + add_599;
assign add_5263 = mulnw_5260 + mulnw_5262;
assign slice_1356 = slice_1352[17:0];
assign addW_6019 = slice_6014 + slice_6011;
assign addW_2112 = slice_2092 + slice_2074;
assign slice_6775 = slice_6774[31:18];
assign slice_2868 = slice_2859[16:8];
assign mulnw_7531 = slice_7529 * slice_7530;
assign subW_3624 = mul_3623 - mul_3615;
assign mul_4380 = slice_4376 * slice_4379;
assign subW_473 = concat_472 - concat_412;
assign slice_5136 = mul_5127[17:0];
assign slice_1229 = slice_1225[17:0];
assign slice_5892 = concat_5779[64:0];
assign slice_1985 = slice_1984[63:32];
assign slice_6648 = slice_6647[32:16];
assign lsl_2741 = mulnw_2740 << 16;
assign mulnw_7404 = slice_7402 * slice_7403;
assign addW_3497 = concat_3491 + subW_3496;
assign concat_4253 = {mul_4248,slice_4252};
assign slice_346 = concat_345[63:32];
assign concat_5009 = {concat_4967,slice_5008};
assign slice_1102 = mul_1093[17:0];
assign slice_5765 = mul_5764[35:18];
assign add_1858 = lsl_1856 + mul_1857;
assign slice_6521 = addW_6435[63:0];
assign mul_2614 = slice_2608 * slice_2610;
assign slice_7277 = addW_7272[17:0];
assign addW_3370 = concat_3081 + subW_3369;
assign slice_4126 = slice_4121[15:0];
assign slice_219 = slice_218[32:16];
assign slice_4882 = slice_4881[31:18];
assign slice_975 = mul_966[17:0];
assign lsl_5638 = mulnw_5637 << 16;
assign mulnw_1731 = slice_1724 * slice_1730;
assign subW_6394 = mul_6393 - mul_6385;
assign lsl_2487 = add_2486 << 8;
assign concat_7150 = {mul_7145,slice_7149};
assign add_3243 = lsl_3241 + mul_3242;
assign slice_3999 = slice_3993[17:0];
assign lsl_92 = mulnw_91 << 16;
assign slice_4755 = slice_4754[32:16];
assign subW_848 = mul_847 - mul_839;
assign addW_5511 = concat_5468 + subW_5510;
assign mulnw_1604 = slice_1603 * slice_1600;
assign subW_6267 = mul_6266 - mul_6258;
assign mul_2360 = slice_2354 * slice_2356;
assign slice_7023 = slice_7016[15:0];
assign mulnw_3116 = slice_3109 * slice_3115;
assign concat_3872 = {addW_3870,slice_3871};
assign mulnw_4628 = slice_4627 * slice_4624;
assign mul_721 = slice_715 * slice_717;
assign addW_5384 = slice_5364 + slice_5344;
assign subW_1477 = mul_1476 - mul_1468;
assign slice_6140 = addW_6139[33:18];
assign subW_2233 = subW_2232 - mul_2226;
assign subW_6896 = subW_6895 - concat_6852;
assign concat_2989 = {concat_2902,slice_2988};
assign concat_3745 = {addW_3743,slice_3744};
assign addW_4501 = slice_4496 + slice_4493;
assign slice_594 = slice_584[7:0];
assign mulnw_5257 = slice_5255 * slice_5256;
assign slice_1350 = addW_1308[31:0];
assign slice_6013 = slice_6008[17:0];
assign slice_2106 = mul_2097[17:0];
assign addW_6769 = concat_6741 + addW_6768;
assign mul_2862 = slice_2859 * slice_2861;
assign slice_7525 = slice_7521[15:0];
assign mul_3618 = slice_3616 * slice_3617;
assign addW_4374 = slice_4287 + slice_4200;
assign add_467 = lsl_465 + mul_466;
assign addW_5130 = slice_5125 + slice_5121;
assign slice_1223 = slice_1222[31:18];
assign addW_5886 = concat_5865 + subW_5885;
assign subW_1979 = subW_1978 - concat_1868;
assign add_6642 = lsl_6633 + add_6641;
assign mul_2735 = slice_2733 * slice_2734;
assign slice_7398 = slice_7394[15:0];
assign concat_3491 = {mul_3486,slice_3490};
assign slice_4247 = slice_4246[31:18];
assign mul_340 = addW_338 * addW_339;
assign add_5003 = lsl_4994 + add_5002;
assign addW_1096 = slice_1091 + slice_1087;
assign addW_5759 = slice_5739 + slice_5699;
assign mulnw_1852 = slice_1851 * slice_1848;
assign addW_6515 = concat_6494 + subW_6514;
assign slice_2608 = slice_2595[7:0];
assign concat_7271 = {concat_7229,slice_7270};
assign subW_3364 = subW_3363 - concat_3253;
assign concat_4120 = {addW_4118,slice_4119};
assign add_4876 = lsl_4867 + add_4875;
assign addW_969 = slice_964 + slice_959;
assign mul_5632 = slice_5626 * slice_5628;
assign slice_1725 = slice_1704[16:8];
assign mul_6388 = slice_6386 * slice_6387;
assign lsl_2481 = mulnw_2480 << 16;
assign slice_7144 = addW_7143[32:16];
assign mulnw_3237 = slice_3236 * slice_3233;
assign slice_3993 = slice_3992[63:32];
assign concat_86 = {mul_80,slice_85};
assign concat_4749 = {addW_4747,slice_4748};
assign mul_842 = slice_840 * slice_841;
assign addW_5505 = add_5491 + add_5504;
assign add_1598 = lsl_1589 + add_1597;
assign mul_6261 = slice_6259 * slice_6260;
assign slice_2354 = slice_2340[7:0];
assign slice_7017 = slice_7016[32:16];
assign slice_3110 = slice_3089[16:8];
assign addW_3866 = slice_3861 + slice_3858;
assign concat_4622 = {mul_4617,slice_4621};
assign slice_715 = slice_702[7:0];
assign subW_5378 = subW_5377 - mul_5371;
assign mul_1471 = slice_1469 * slice_1470;
assign concat_6134 = {addW_6132,slice_6133};
assign slice_2227 = mul_2226[35:18];
assign add_6890 = lsl_6881 + add_6889;
assign subW_2983 = concat_2982 - concat_2922;
assign addW_3739 = slice_3734 + slice_3731;
assign slice_4495 = slice_4488[17:0];
assign slice_588 = slice_577[16:8];
assign lsl_5251 = add_5250 << 8;
assign add_1344 = lsl_1342 + mul_1343;
assign concat_6007 = {addW_6005,slice_6006};
assign addW_2100 = slice_2095 + slice_2091;
assign add_6763 = mulnw_6760 + mulnw_6762;
assign slice_2856 = concat_2855[63:32];
assign slice_7519 = addW_7477[32:0];
assign slice_3612 = addW_3611[33:18];
assign subW_4368 = subW_4367 - concat_4324;
assign mulnw_461 = slice_460 * slice_457;
assign mul_5124 = slice_5121 * slice_5123;
assign subW_1217 = subW_1216 - concat_1173;
assign subW_5880 = subW_5879 - mul_5873;
assign subW_1973 = concat_1972 - concat_1912;
assign slice_6636 = slice_6610[7:0];
assign addW_2729 = slice_2642 + slice_2557;
assign slice_7392 = slice_7391[32:16];
assign slice_3485 = slice_3484[31:18];
assign addW_4241 = concat_4213 + addW_4240;
assign slice_334 = slice_330[17:0];
assign slice_4997 = slice_4971[7:0];
assign mul_1090 = slice_1087 * slice_1089;
assign slice_5753 = mul_5744[17:0];
assign add_1846 = lsl_1837 + add_1845;
assign subW_6509 = subW_6508 - mul_6502;
assign slice_2602 = mul_2601[31:16];
assign add_7265 = lsl_7256 + add_7264;
assign subW_3358 = concat_3357 - concat_3297;
assign mul_4114 = slice_4108 * slice_4110;
assign addW_207 = concat_164 + subW_206;
assign slice_4870 = slice_4844[7:0];
assign mul_963 = slice_959 * slice_962;
assign slice_5626 = slice_5611[7:0];
assign add_1719 = mulnw_1716 + mulnw_1718;
assign slice_6382 = slice_6381[31:18];
assign mul_2475 = slice_2473 * slice_2474;
assign concat_7138 = {addW_7136,slice_7137};
assign add_3231 = lsl_3222 + add_3230;
assign subW_3987 = concat_3986 - concat_3948;
assign mul_80 = slice_77 * slice_79;
assign slice_4743 = concat_4719[31:0];
assign slice_836 = addW_835[33:18];
assign mulnw_5499 = slice_5492 * slice_5498;
assign slice_1592 = slice_1582[7:0];
assign slice_6255 = slice_6169[63:0];
assign slice_2348 = mul_2347[31:16];
assign addW_7011 = concat_6901 + subW_7010;
assign add_3104 = mulnw_3101 + mulnw_3103;
assign slice_3860 = slice_3855[17:0];
assign slice_4616 = addW_4615[32:16];
assign slice_709 = mul_708[31:16];
assign slice_5372 = mul_5371[35:18];
assign slice_1465 = addW_1464[33:18];
assign addW_6128 = slice_6123 + slice_6120;
assign addW_2221 = slice_2201 + slice_2161;
assign slice_6884 = slice_6858[7:0];
assign add_2977 = lsl_2975 + mul_2976;
assign slice_3733 = slice_3727[17:0];
assign slice_4489 = slice_4488[31:18];
assign mul_582 = slice_577 * slice_581;
assign lsl_5245 = mulnw_5244 << 16;
assign mulnw_1338 = slice_1337 * slice_1334;
assign addW_6001 = slice_5996 + slice_5993;
assign mul_2094 = slice_2091 * slice_2093;
assign mulnw_6757 = slice_6755 * slice_6756;
assign mul_2850 = addW_2848 * addW_2849;
assign add_7513 = lsl_7511 + mul_7512;
assign addW_3606 = concat_3600 + subW_3605;
assign add_4362 = lsl_4353 + add_4361;
assign add_455 = lsl_446 + add_454;
assign slice_5118 = concat_5117[63:32];
assign add_1211 = lsl_1202 + add_1210;
assign slice_5874 = mul_5873[35:18];
assign mul_1967 = addW_1965 * addW_1966;
assign slice_6630 = slice_6612[15:8];
assign concat_2723 = {addW_2721,slice_2722};
assign subW_7386 = subW_7385 - concat_7364;
assign addW_3479 = concat_3473 + subW_3478;
assign add_4235 = mulnw_4232 + mulnw_4234;
assign slice_328 = slice_307[31:0];
assign slice_4991 = slice_4973[15:8];
assign slice_1084 = mul_1053[15:0];
assign addW_5747 = slice_5742 + slice_5738;
assign slice_1840 = slice_1830[7:0];
assign slice_6503 = mul_6502[35:18];
assign addW_2596 = slice_2576 + slice_2558;
assign slice_7259 = slice_7233[7:0];
assign mul_3352 = addW_3350 * addW_3351;
assign slice_4108 = slice_4086[7:0];
assign addW_201 = add_187 + add_200;
assign slice_4864 = slice_4846[15:8];
assign slice_957 = slice_869[63:0];
assign slice_5620 = mul_5619[31:16];
assign mulnw_1713 = slice_1711 * slice_1712;
assign add_6376 = lsl_6367 + add_6375;
assign slice_2469 = slice_2468[32:16];
assign addW_7132 = slice_7127 + slice_7124;
assign slice_3225 = slice_3215[7:0];
assign mul_3981 = addW_3979 * addW_3980;
assign addW_4737 = concat_4731 + subW_4736;
assign slice_830 = mul_799[15:0];
assign slice_5493 = slice_5472[16:8];
assign slice_1586 = slice_1576[16:8];
assign addW_6249 = concat_6206 + subW_6248;
assign slice_2342 = slice_2341[64:32];
assign subW_7005 = subW_7004 - concat_6983;
assign mulnw_3098 = slice_3096 * slice_3097;
assign concat_3854 = {addW_3852,slice_3853};
assign concat_4610 = {addW_4608,slice_4609};
assign addW_703 = slice_683 + slice_665;
assign slice_5366 = slice_5347[31:0];
assign addW_1459 = concat_1453 + subW_1458;
assign slice_6122 = slice_6117[17:0];
assign slice_2215 = mul_2206[17:0];
assign slice_6878 = slice_6860[15:8];
assign mulnw_2971 = slice_2970 * slice_2967;
assign slice_3727 = slice_3726[63:32];
assign addW_4483 = concat_4373 + subW_4482;
assign slice_576 = slice_575[64:32];
assign mul_5239 = slice_5237 * slice_5238;
assign add_1332 = lsl_1323 + add_1331;
assign slice_5995 = slice_5989[17:0];
assign slice_2088 = mul_2079[17:0];
assign lsl_6751 = add_6750 << 8;
assign slice_2844 = slice_2840[17:0];
assign mulnw_7507 = slice_7506 * slice_7503;
assign concat_3600 = {mul_3595,slice_3599};
assign slice_4356 = slice_4330[7:0];
assign slice_449 = slice_439[7:0];
assign mul_5112 = addW_5110 * addW_5111;
assign slice_1205 = slice_1179[7:0];
assign addW_5868 = slice_5826 + slice_5786;
assign slice_1961 = addW_1957[17:0];
assign mulnw_6624 = slice_6617 * slice_6623;
assign slice_2717 = mul_2686[15:0];
assign subW_7380 = mul_7379 - mul_7371;
assign concat_3473 = {mul_3468,slice_3472};
assign mulnw_4229 = slice_4227 * slice_4228;
assign mul_322 = addW_320 * addW_321;
assign mulnw_4985 = slice_4978 * slice_4984;
assign lsl_1078 = add_1077 << 8;
assign mul_5741 = slice_5738 * slice_5740;
assign slice_1834 = slice_1825[16:8];
assign addW_6497 = slice_6477 + slice_6437;
assign slice_2590 = mul_2581[17:0];
assign slice_7253 = slice_7235[15:8];
assign slice_3346 = addW_3342[17:0];
assign add_4102 = lsl_4100 + mul_4101;
assign mulnw_195 = slice_188 * slice_194;
assign mulnw_4858 = slice_4851 * slice_4857;
assign concat_951 = {addW_949,slice_950};
assign slice_5614 = slice_5613[64:32];
assign slice_1707 = slice_1703[15:0];
assign slice_6370 = slice_6344[7:0];
assign add_2463 = lsl_2454 + add_2462;
assign slice_7126 = slice_7121[17:0];
assign slice_3219 = slice_3210[16:8];
assign slice_3975 = addW_3971[17:0];
assign slice_68 = mul_59[17:0];
assign concat_4731 = {mul_4726,slice_4730};
assign lsl_824 = add_823 << 8;
assign add_5487 = mulnw_5484 + mulnw_5486;
assign mul_1580 = slice_1576 * slice_1579;
assign addW_6243 = add_6229 + add_6242;
assign slice_2336 = concat_2312[31:0];
assign subW_6999 = mul_6998 - mul_6990;
assign slice_3092 = slice_3088[15:0];
assign mul_3848 = slice_3842 * slice_3844;
assign addW_4604 = slice_4599 + slice_4596;
assign slice_697 = mul_688[17:0];
assign subW_5360 = subW_5359 - mul_5353;
assign concat_1453 = {mul_1448,slice_1452};
assign concat_6116 = {addW_6114,slice_6115};
assign addW_2209 = slice_2204 + slice_2200;
assign mulnw_6872 = slice_6865 * slice_6871;
assign add_2965 = lsl_2956 + add_2964;
assign subW_3721 = concat_3720 - concat_3660;
assign subW_4477 = subW_4476 - concat_4455;
assign slice_570 = concat_569[255:128];
assign addW_5233 = slice_5146 + slice_5061;
assign slice_1326 = slice_1316[7:0];
assign slice_5989 = slice_5988[63:32];
assign addW_2082 = slice_2077 + slice_2072;
assign lsl_6745 = mulnw_6744 << 16;
assign slice_2838 = slice_2817[31:0];
assign add_7501 = lsl_7492 + add_7500;
assign slice_3594 = slice_3593[31:18];
assign slice_4350 = slice_4332[15:8];
assign slice_443 = slice_434[16:8];
assign slice_5106 = slice_5102[17:0];
assign slice_1199 = slice_1181[15:8];
assign slice_5862 = mul_5831[15:0];
assign addW_1955 = slice_1913 + slice_1872;
assign slice_6618 = slice_6613[15:8];
assign lsl_2711 = add_2710 << 8;
assign mul_7374 = slice_7372 * slice_7373;
assign slice_3467 = slice_3466[31:18];
assign lsl_4223 = add_4222 << 8;
assign slice_316 = slice_312[17:0];
assign slice_4979 = slice_4974[15:8];
assign lsl_1072 = mulnw_1071 << 16;
assign slice_5735 = mul_5704[15:0];
assign mul_1828 = slice_1825 * slice_1827;
assign slice_6491 = mul_6482[17:0];
assign addW_2584 = slice_2579 + slice_2575;
assign mulnw_7247 = slice_7240 * slice_7246;
assign addW_3340 = slice_3298 + slice_3257;
assign mulnw_4096 = slice_4095 * slice_4092;
assign slice_189 = slice_168[16:8];
assign slice_4852 = slice_4847[15:8];
assign mul_945 = slice_939 * slice_941;
assign addW_5608 = slice_5342 + slice_5054;
assign slice_1701 = addW_1700[256:128];
assign slice_6364 = slice_6346[15:8];
assign slice_2457 = slice_2431[7:0];
assign concat_7120 = {addW_7118,slice_7119};
assign mul_3213 = slice_3210 * slice_3212;
assign addW_3969 = slice_3949 + slice_3907;
assign addW_62 = slice_57 + slice_53;
assign slice_4725 = addW_4724[33:18];
assign lsl_818 = mulnw_817 << 16;
assign mulnw_5481 = slice_5479 * slice_5480;
assign addW_1574 = slice_1487 + slice_1401;
assign mulnw_6237 = slice_6230 * slice_6236;
assign addW_2330 = concat_2324 + subW_2329;
assign mul_6993 = slice_6991 * slice_6992;
assign addW_3086 = slice_2820 + slice_2556;
assign slice_3842 = slice_3820[7:0];
assign slice_4598 = slice_4593[17:0];
assign addW_691 = slice_686 + slice_682;
assign slice_5354 = mul_5353[35:18];
assign slice_1447 = slice_1446[31:18];
assign mul_6110 = slice_6104 * slice_6106;
assign mul_2203 = slice_2200 * slice_2202;
assign slice_6866 = slice_6861[15:8];
assign slice_2959 = slice_2949[7:0];
assign add_3715 = lsl_3713 + mul_3714;
assign subW_4471 = mul_4470 - mul_4462;
assign concat_564 = {addW_562,slice_563};
assign concat_5227 = {addW_5225,slice_5226};
assign slice_1320 = slice_1310[16:8];
assign subW_5983 = concat_5982 - concat_5922;
assign mul_2076 = slice_2072 * slice_2075;
assign mul_6739 = slice_6737 * slice_6738;
assign mul_2832 = addW_2830 * addW_2831;
assign slice_7495 = slice_7485[7:0];
assign addW_3588 = concat_3560 + addW_3587;
assign mulnw_4344 = slice_4337 * slice_4343;
assign mul_437 = slice_434 * slice_436;
assign slice_5100 = slice_5055[31:0];
assign mulnw_1193 = slice_1186 * slice_1192;
assign lsl_5856 = add_5855 << 8;
assign addW_1949 = add_1935 + add_1948;
assign slice_6612 = slice_6606[15:0];
assign lsl_2705 = mulnw_2704 << 16;
assign slice_7368 = addW_7367[33:18];
assign concat_3461 = {addW_3459,slice_3460};
assign lsl_4217 = mulnw_4216 << 16;
assign slice_310 = slice_28[127:0];
assign slice_4973 = slice_4968[15:0];
assign mul_1066 = slice_1060 * slice_1062;
assign lsl_5729 = add_5728 << 8;
assign slice_1822 = concat_1821[63:32];
assign addW_6485 = slice_6480 + slice_6476;
assign mul_2578 = slice_2575 * slice_2577;
assign slice_7241 = slice_7236[15:8];
assign addW_3334 = add_3320 + add_3333;
assign concat_4090 = {mul_4085,slice_4089};
assign add_183 = mulnw_180 + mulnw_182;
assign slice_4846 = slice_4840[15:0];
assign slice_939 = slice_917[7:0];
assign subW_5602 = subW_5601 - concat_5513;
assign addW_1695 = slice_868 + slice_13;
assign mulnw_6358 = slice_6351 * slice_6357;
assign slice_2451 = slice_2433[15:8];
assign addW_7114 = slice_7109 + slice_7106;
assign slice_3207 = concat_3206[63:32];
assign subW_3963 = subW_3962 - mul_3956;
assign mul_56 = slice_53 * slice_55;
assign concat_4719 = {addW_4717,slice_4718};
assign mul_812 = slice_806 * slice_808;
assign slice_5475 = addW_5471[15:0];
assign subW_1568 = subW_1567 - concat_1524;
assign slice_6231 = slice_6210[16:8];
assign concat_2324 = {mul_2319,slice_2323};
assign slice_6987 = addW_6986[33:18];
assign slice_3080 = concat_3079[255:128];
assign add_3836 = lsl_3834 + mul_3835;
assign concat_4592 = {addW_4590,slice_4591};
assign mul_685 = slice_682 * slice_684;
assign slice_5348 = slice_5347[63:32];
assign addW_1441 = concat_1413 + addW_1440;
assign slice_6104 = slice_6082[7:0];
assign slice_2197 = mul_2166[15:0];
assign slice_6860 = addW_6855[15:0];
assign slice_2953 = slice_2944[16:8];
assign mulnw_3709 = slice_3708 * slice_3705;
assign mul_4465 = slice_4463 * slice_4464;
assign slice_558 = mul_549[17:0];
assign slice_5221 = mul_5190[15:0];
assign mul_1314 = slice_1310 * slice_1313;
assign add_5977 = lsl_5975 + mul_5976;
assign slice_2070 = slice_1983[63:0];
assign slice_6733 = slice_6732[128:64];
assign slice_2826 = slice_2822[17:0];
assign slice_7489 = slice_7479[16:8];
assign add_3582 = mulnw_3579 + mulnw_3581;
assign slice_4338 = slice_4333[15:8];
assign slice_431 = concat_430[63:32];
assign add_5094 = lsl_5092 + mul_5093;
assign slice_1187 = slice_1182[15:8];
assign lsl_5850 = mulnw_5849 << 16;
assign mulnw_1943 = slice_1936 * slice_1942;
assign slice_6606 = addW_6605[65:33];
assign mul_2699 = slice_2693 * slice_2695;
assign addW_7362 = concat_7356 + subW_7361;
assign slice_3455 = mul_3424[15:0];
assign mul_4211 = slice_4209 * slice_4210;
assign slice_304 = concat_209[63:0];
assign concat_4967 = {addW_4965,slice_4966};
assign slice_1060 = slice_1046[7:0];
assign lsl_5723 = mulnw_5722 << 16;
assign mul_1816 = addW_1814 * addW_1815;
assign mul_6479 = slice_6476 * slice_6478;
assign slice_2572 = mul_2563[17:0];
assign slice_7235 = slice_7230[15:0];
assign mulnw_3328 = slice_3321 * slice_3327;
assign slice_4084 = slice_4083[32:16];
assign mulnw_177 = slice_175 * slice_176;
assign slice_4840 = slice_4839[64:32];
assign add_933 = lsl_931 + mul_932;
assign subW_5596 = concat_5595 - concat_5557;
assign slice_1689 = concat_1397[127:0];
assign slice_6352 = slice_6347[15:8];
assign mulnw_2445 = slice_2438 * slice_2444;
assign slice_7108 = slice_7102[17:0];
assign mul_3201 = addW_3199 * addW_3200;
assign slice_3957 = mul_3956[35:18];
assign slice_50 = mul_38[17:0];
assign addW_4713 = slice_4708 + slice_4705;
assign slice_806 = slice_793[7:0];
assign addW_5469 = slice_5449 + slice_5430;
assign add_1562 = lsl_1553 + add_1561;
assign add_6225 = mulnw_6222 + mulnw_6224;
assign slice_2318 = addW_2317[33:18];
assign addW_6981 = concat_6953 + addW_6980;
assign concat_3074 = {addW_3072,slice_3073};
assign mulnw_3830 = slice_3829 * slice_3826;
assign addW_4586 = slice_4581 + slice_4578;
assign slice_679 = mul_670[17:0];
assign slice_5342 = slice_5053[127:0];
assign add_1435 = mulnw_1432 + mulnw_1434;
assign add_6098 = lsl_6096 + mul_6097;
assign lsl_2191 = add_2190 << 8;
assign concat_6854 = {concat_6834,slice_6853};
assign mul_2947 = slice_2944 * slice_2946;
assign add_3703 = lsl_3694 + add_3702;
assign slice_4459 = addW_4458[33:18];
assign addW_552 = slice_547 + slice_543;
assign lsl_5215 = add_5214 << 8;
assign addW_1308 = slice_1221 + slice_1135;
assign mulnw_5971 = slice_5970 * slice_5967;
assign concat_2064 = {addW_2062,slice_2063};
assign slice_6727 = addW_6726[257:129];
assign slice_2820 = slice_2555[127:0];
assign mul_7483 = slice_7479 * slice_7482;
assign mulnw_3576 = slice_3574 * slice_3575;
assign slice_4332 = addW_4327[15:0];
assign mul_425 = addW_423 * addW_424;
assign mulnw_5088 = slice_5087 * slice_5084;
assign slice_1181 = addW_1176[15:0];
assign mul_5844 = slice_5838 * slice_5840;
assign slice_1937 = slice_1916[16:8];
assign addW_6600 = concat_6557 + subW_6599;
assign slice_2693 = slice_2680[7:0];
assign concat_7356 = {mul_7351,slice_7355};
assign lsl_3449 = add_3448 << 8;
assign slice_4205 = slice_4204[128:64];
assign addW_298 = concat_275 + subW_297;
assign mul_4961 = slice_4955 * slice_4957;
assign slice_1054 = mul_1053[31:16];
assign mul_5717 = slice_5711 * slice_5713;
assign slice_1810 = slice_1806[17:0];
assign slice_6473 = mul_6442[15:0];
assign addW_2566 = slice_2561 + slice_2553;
assign concat_7229 = {addW_7227,slice_7228};
assign slice_3322 = slice_3301[16:8];
assign concat_4078 = {concat_3991,slice_4077};
assign slice_171 = addW_167[15:0];
assign subW_4834 = concat_4833 - concat_4795;
assign mulnw_927 = slice_926 * slice_923;
assign mul_5590 = addW_5588 * addW_5589;
assign addW_1683 = concat_1573 + subW_1682;
assign slice_6346 = slice_6340[15:0];
assign slice_2439 = slice_2434[15:8];
assign slice_7102 = slice_7101[63:32];
assign slice_3195 = slice_3191[17:0];
assign slice_3951 = slice_3910[31:0];
assign addW_44 = slice_36 + slice_25;
assign slice_4707 = slice_4702[17:0];
assign slice_800 = mul_799[31:16];
assign subW_5463 = subW_5462 - mul_5456;
assign slice_1556 = slice_1530[7:0];
assign mulnw_6219 = slice_6217 * slice_6218;
assign concat_2312 = {addW_2310,slice_2311};
assign add_6975 = mulnw_6972 + mulnw_6974;
assign slice_3068 = mul_3059[17:0];
assign concat_3824 = {mul_3819,slice_3823};
assign slice_4580 = slice_4574[17:0];
assign addW_673 = slice_668 + slice_663;
assign concat_5336 = {addW_5334,slice_5335};
assign mulnw_1429 = slice_1427 * slice_1428;
assign mulnw_6092 = slice_6091 * slice_6088;
assign lsl_2185 = mulnw_2184 << 16;
assign subW_6848 = mul_6847 - mul_6839;
assign slice_2941 = concat_2940[63:32];
assign slice_3697 = slice_3687[7:0];
assign addW_4453 = concat_4425 + addW_4452;
assign mul_546 = slice_543 * slice_545;
assign lsl_5209 = mulnw_5208 << 16;
assign subW_1302 = subW_1301 - concat_1258;
assign add_5965 = lsl_5956 + add_5964;
assign mul_2058 = slice_2052 * slice_2054;
assign concat_6721 = {addW_6719,slice_6720};
assign slice_2814 = concat_2723[63:0];
assign addW_7477 = slice_7390 + slice_7304;
assign lsl_3570 = add_3569 << 8;
assign concat_4326 = {concat_4306,slice_4325};
assign slice_419 = slice_415[17:0];
assign add_5082 = lsl_5073 + add_5081;
assign concat_1175 = {concat_1155,slice_1174};
assign slice_5838 = slice_5825[7:0];
assign add_1931 = mulnw_1928 + mulnw_1930;
assign addW_6594 = add_6580 + add_6593;
assign slice_2687 = mul_2686[31:16];
assign slice_7350 = slice_7349[31:18];
assign lsl_3443 = mulnw_3442 << 16;
assign slice_4199 = addW_4198[256:128];
assign subW_292 = subW_291 - mul_285;
assign slice_4955 = slice_4933[7:0];
assign slice_1048 = addW_1047[64:32];
assign slice_5711 = slice_5697[7:0];
assign slice_1804 = slice_1784[31:0];
assign lsl_6467 = add_6466 << 8;
assign mul_2560 = slice_2553 * slice_2559;
assign mul_7223 = slice_7217 * slice_7219;
assign add_3316 = mulnw_3313 + mulnw_3315;
assign subW_4072 = concat_4071 - concat_4011;
assign addW_165 = slice_145 + slice_126;
assign mul_4828 = addW_4826 * addW_4827;
assign concat_921 = {mul_916,slice_920};
assign slice_5584 = addW_5580[17:0];
assign subW_1677 = subW_1676 - concat_1655;
assign slice_6340 = addW_6339[64:32];
assign slice_2433 = slice_2427[15:0];
assign subW_7096 = concat_7095 - concat_7057;
assign slice_3189 = slice_3169[31:0];
assign addW_3945 = add_3931 + add_3944;
assign mul_38 = slice_36 * slice_37;
assign concat_4701 = {addW_4699,slice_4700};
assign slice_794 = addW_753[32:0];
assign slice_5457 = mul_5456[35:18];
assign slice_1550 = slice_1532[15:8];
assign slice_6213 = addW_6209[15:0];
assign addW_2306 = slice_2301 + slice_2298;
assign mulnw_6969 = slice_6967 * slice_6968;
assign addW_3062 = slice_3057 + slice_3053;
assign slice_3818 = slice_3817[32:16];
assign slice_4574 = slice_4573[63:32];
assign mul_667 = slice_663 * slice_666;
assign slice_5330 = mul_5321[17:0];
assign lsl_1423 = add_1422 << 8;
assign concat_6086 = {mul_6081,slice_6085};
assign mul_2179 = slice_2173 * slice_2175;
assign mul_6842 = slice_6840 * slice_6841;
assign mul_2935 = addW_2933 * addW_2934;
assign concat_7598 = {addW_7596,slice_7597};
assign slice_3691 = slice_3682[16:8];
assign add_4447 = mulnw_4444 + mulnw_4446;
assign slice_540 = concat_539[63:32];
assign mul_5203 = slice_5197 * slice_5199;
assign add_1296 = lsl_1287 + add_1295;
assign slice_5959 = slice_5949[7:0];
assign slice_2052 = slice_2030[7:0];
assign slice_6715 = concat_6602[63:0];
assign addW_2808 = concat_2787 + subW_2807;
assign subW_7471 = subW_7470 - concat_7449;
assign lsl_3564 = mulnw_3563 << 16;
assign subW_4320 = mul_4319 - mul_4311;
assign slice_413 = slice_393[31:0];
assign slice_5076 = slice_5066[7:0];
assign subW_1169 = mul_1168 - mul_1160;
assign slice_5832 = mul_5831[31:16];
assign mulnw_1925 = slice_1923 * slice_1924;
assign mulnw_6588 = slice_6581 * slice_6587;
assign addW_2681 = slice_2661 + slice_2643;
assign addW_7344 = concat_7316 + addW_7343;
assign mul_3437 = slice_3431 * slice_3433;
assign addW_4193 = concat_3904 + subW_4192;
assign slice_286 = mul_285[35:18];
assign add_4949 = lsl_4947 + mul_4948;
assign slice_1042 = concat_1041[127:64];
assign slice_5705 = mul_5704[31:16];
assign mul_1798 = addW_1796 * addW_1797;
assign lsl_6461 = mulnw_6460 << 16;
assign slice_2554 = IN2[511:0];
assign slice_7217 = slice_7195[7:0];
assign mulnw_3310 = slice_3308 * slice_3309;
assign add_4066 = lsl_4064 + mul_4065;
assign subW_159 = subW_158 - mul_152;
assign slice_4822 = addW_4818[17:0];
assign slice_915 = addW_914[32:16];
assign addW_5578 = slice_5558 + slice_5517;
assign subW_1671 = mul_1670 - mul_1662;
assign addW_6334 = concat_6291 + subW_6333;
assign slice_2427 = addW_2426[65:33];
assign mul_7090 = addW_7088 * addW_7089;
assign mul_3183 = addW_3181 * addW_3182;
assign mulnw_3939 = slice_3932 * slice_3938;
assign slice_32 = slice_31[31:18];
assign mul_4695 = slice_4689 * slice_4691;
assign addW_788 = add_774 + add_787;
assign slice_5451 = slice_5432[31:0];
assign mulnw_1544 = slice_1537 * slice_1543;
assign addW_6207 = slice_6187 + slice_6167;
assign slice_2300 = slice_2295[17:0];
assign lsl_6963 = add_6962 << 8;
assign mul_3056 = slice_3053 * slice_3055;
assign concat_3812 = {concat_3725,slice_3811};
assign subW_4568 = concat_4567 - concat_4507;
assign slice_661 = addW_574[63:0];
assign addW_5324 = slice_5319 + slice_5315;
assign lsl_1417 = mulnw_1416 << 16;
assign slice_6080 = slice_6079[32:16];
assign slice_2173 = slice_2159[7:0];
assign slice_6836 = slice_6835[31:18];
assign slice_2929 = slice_2925[17:0];
assign slice_7592 = concat_7299[128:0];
assign mul_3685 = slice_3682 * slice_3684;
assign mulnw_4441 = slice_4439 * slice_4440;
assign mul_534 = addW_532 * addW_533;
assign slice_5197 = slice_5184[7:0];
assign slice_1290 = slice_1264[7:0];
assign slice_5953 = slice_5944[16:8];
assign add_2046 = lsl_2044 + mul_2045;
assign addW_6709 = concat_6688 + subW_6708;
assign subW_2802 = subW_2801 - mul_2795;
assign subW_7465 = mul_7464 - mul_7456;
assign mul_3558 = slice_3556 * slice_3557;
assign mul_4314 = slice_4312 * slice_4313;
assign mul_407 = addW_405 * addW_406;
assign slice_5070 = slice_5057[16:8];
assign mul_1163 = slice_1161 * slice_1162;
assign slice_5826 = addW_5785[32:0];
assign slice_1919 = slice_1915[15:0];
assign slice_6582 = slice_6561[16:8];
assign slice_2675 = mul_2666[17:0];
assign add_7338 = mulnw_7335 + mulnw_7337;
assign slice_3431 = slice_3418[7:0];
assign subW_4187 = subW_4186 - concat_4076;
assign addW_280 = slice_258 + slice_218;
assign mulnw_4943 = slice_4942 * slice_4939;
assign concat_1036 = {addW_1034,slice_1035};
assign slice_5699 = slice_5698[64:32];
assign slice_1792 = slice_1788[17:0];
assign mul_6455 = slice_6449 * slice_6451;
assign slice_2548 = IN1[511:0];
assign add_7211 = lsl_7209 + mul_7210;
assign slice_3304 = slice_3300[15:0];
assign mulnw_4060 = slice_4059 * slice_4056;
assign slice_153 = mul_152[35:18];
assign addW_4816 = slice_4796 + slice_4754;
assign concat_909 = {addW_907,slice_908};
assign subW_5572 = subW_5571 - mul_5565;
assign mul_1665 = slice_1663 * slice_1664;
assign addW_6328 = add_6314 + add_6327;
assign slice_2421 = concat_2397[31:0];
assign slice_7084 = addW_7080[17:0];
assign slice_3177 = slice_3173[17:0];
assign slice_3933 = slice_3912[16:8];
assign slice_4689 = slice_4667[7:0];
assign mulnw_782 = slice_775 * slice_781;
assign subW_5445 = subW_5444 - mul_5438;
assign slice_1538 = slice_1533[15:8];
assign subW_6201 = subW_6200 - mul_6194;
assign concat_2294 = {addW_2292,slice_2293};
assign lsl_6957 = mulnw_6956 << 16;
assign slice_3050 = concat_3049[63:32];
assign subW_3806 = concat_3805 - concat_3745;
assign add_4562 = lsl_4560 + mul_4561;
assign concat_655 = {addW_653,slice_654};
assign mul_5318 = slice_5315 * slice_5317;
assign mul_1411 = slice_1409 * slice_1410;
assign concat_6074 = {concat_5987,slice_6073};
assign slice_2167 = mul_2166[31:16];
assign subW_6830 = mul_6829 - mul_6821;
assign slice_2923 = slice_2903[31:0];
assign addW_7586 = concat_7476 + subW_7585;
assign slice_3679 = concat_3678[63:32];
assign lsl_4435 = add_4434 << 8;
assign slice_528 = slice_524[17:0];
assign slice_5191 = mul_5190[31:16];
assign slice_1284 = slice_1266[15:8];
assign mul_5947 = slice_5944 * slice_5946;
assign mulnw_2040 = slice_2039 * slice_2036;
assign subW_6703 = subW_6702 - mul_6696;
assign slice_2796 = mul_2795[35:18];
assign mul_7459 = slice_7457 * slice_7458;
assign addW_3552 = slice_3465 + slice_3380;
assign slice_4308 = slice_4307[31:18];
assign slice_401 = slice_397[17:0];
assign mul_5064 = slice_5057 * slice_5063;
assign slice_1157 = slice_1156[31:18];
assign addW_5820 = add_5806 + add_5819;
assign slice_1913 = addW_1871[32:0];
assign add_6576 = mulnw_6573 + mulnw_6575;
assign addW_2669 = slice_2664 + slice_2660;
assign mulnw_7332 = slice_7330 * slice_7331;
assign slice_3425 = mul_3424[31:16];
assign subW_4181 = concat_4180 - concat_4120;
assign slice_274 = concat_273[63:32];
assign concat_4937 = {mul_4932,slice_4936};
assign mul_1030 = slice_1024 * slice_1026;
assign slice_5693 = concat_5669[31:0];
assign slice_1786 = slice_1785[31:18];
assign slice_6449 = slice_6434[7:0];
assign concat_2542 = {addW_2540,slice_2541};
assign mulnw_7205 = slice_7204 * slice_7201;
assign slice_3298 = addW_3256[32:0];
assign add_4054 = lsl_4045 + add_4053;
assign slice_147 = slice_128[31:0];
assign subW_4810 = subW_4809 - mul_4803;
assign addW_903 = slice_898 + slice_895;
assign slice_5566 = mul_5565[35:18];
assign slice_1659 = addW_1658[33:18];
assign mulnw_6322 = slice_6315 * slice_6321;
assign addW_2415 = concat_2409 + subW_2414;
assign addW_7078 = slice_7058 + slice_7016;
assign slice_3171 = slice_3170[31:18];
assign add_3927 = mulnw_3924 + mulnw_3926;
assign add_4683 = lsl_4681 + mul_4682;
assign slice_776 = slice_755[16:8];
assign slice_5439 = mul_5438[35:18];
assign slice_1532 = addW_1527[15:0];
assign slice_6195 = mul_6194[35:18];
assign mul_2288 = slice_2282 * slice_2284;
assign mul_6951 = slice_6949 * slice_6950;
assign mul_3044 = addW_3042 * addW_3043;
assign add_3800 = lsl_3798 + mul_3799;
assign mulnw_4556 = slice_4555 * slice_4552;
assign addW_649 = slice_644 + slice_641;
assign slice_5312 = concat_5311[65:33];
assign slice_1405 = addW_1404[128:64];
assign subW_6068 = concat_6067 - concat_6007;
assign slice_2161 = addW_2160[64:32];
assign mul_6824 = slice_6822 * slice_6823;
assign mul_2917 = addW_2915 * addW_2916;
assign subW_7580 = subW_7579 - concat_7558;
assign mul_3673 = addW_3671 * addW_3672;
assign lsl_4429 = mulnw_4428 << 16;
assign slice_522 = addW_480[31:0];
assign addW_5185 = slice_5165 + slice_5147;
assign mulnw_1278 = slice_1271 * slice_1277;
assign slice_5941 = concat_5940[63:32];
assign concat_2034 = {mul_2029,slice_2033};
assign slice_6697 = mul_6696[35:18];
assign addW_2790 = slice_2770 + slice_2730;
assign slice_7453 = addW_7452[33:18];
assign concat_3546 = {addW_3544,slice_3545};
assign subW_4302 = mul_4301 - mul_4293;
assign slice_395 = slice_394[31:18];
assign addW_5058 = slice_2554 + slice_27;
assign subW_1151 = mul_1150 - mul_1142;
assign mulnw_5814 = slice_5807 * slice_5813;
assign add_1907 = lsl_1905 + mul_1906;
assign mulnw_6570 = slice_6568 * slice_6569;
assign mul_2663 = slice_2660 * slice_2662;
assign lsl_7326 = add_7325 << 8;
assign addW_3419 = slice_3399 + slice_3381;
assign mul_4175 = addW_4173 * addW_4174;
assign mul_268 = addW_266 * addW_267;
assign slice_4931 = slice_4930[32:16];
assign slice_1024 = slice_1002[7:0];
assign addW_5687 = concat_5681 + subW_5686;
assign subW_1780 = subW_1779 - concat_1758;
assign slice_6443 = mul_6442[31:16];
assign slice_2536 = concat_2422[64:0];
assign concat_7199 = {mul_7194,slice_7198};
assign add_3292 = lsl_3290 + mul_3291;
assign slice_4048 = slice_4038[7:0];
assign subW_141 = subW_140 - mul_134;
assign slice_4804 = mul_4803[35:18];
assign slice_897 = slice_892[17:0];
assign slice_5560 = addW_5519[31:0];
assign addW_1653 = concat_1625 + addW_1652;
assign slice_6316 = slice_6295[16:8];
assign concat_2409 = {mul_2404,slice_2408};
assign subW_7072 = subW_7071 - mul_7065;
assign subW_3165 = subW_3164 - concat_3143;
assign mulnw_3921 = slice_3919 * slice_3920;
assign mulnw_4677 = slice_4676 * slice_4673;
assign add_770 = mulnw_767 + mulnw_769;
assign slice_5433 = slice_5432[63:32];
assign concat_1526 = {concat_1506,slice_1525};
assign slice_6189 = slice_6170[31:0];
assign slice_2282 = slice_2260[7:0];
assign slice_6945 = slice_6944[32:16];
assign slice_3038 = slice_3034[17:0];
assign mulnw_3794 = slice_3793 * slice_3790;
assign add_4550 = lsl_4541 + add_4549;
assign slice_643 = addW_638[17:0];
assign add_5306 = lsl_5304 + mul_5305;
assign concat_1399 = {concat_1133,slice_1398};
assign add_6062 = lsl_6060 + mul_6061;
assign slice_2155 = concat_2154[127:64];
assign slice_6818 = slice_6732[63:0];
assign slice_2911 = slice_2907[17:0];
assign subW_7574 = mul_7573 - mul_7565;
assign slice_3667 = slice_3663[17:0];
assign mul_4423 = slice_4421 * slice_4422;
assign add_516 = lsl_514 + mul_515;
assign slice_5179 = mul_5170[17:0];
assign slice_1272 = slice_1267[15:8];
assign mul_5935 = addW_5933 * addW_5934;
assign slice_2028 = addW_2027[32:16];
assign addW_6691 = slice_6649 + slice_6609;
assign slice_2784 = mul_2775[17:0];
assign addW_7447 = concat_7441 + subW_7446;
assign slice_3540 = mul_3509[15:0];
assign mul_4296 = slice_4294 * slice_4295;
assign subW_389 = subW_388 - concat_345;
assign addW_5052 = slice_2548 + slice_10;
assign mul_1145 = slice_1143 * slice_1144;
assign slice_5808 = slice_5787[16:8];
assign mulnw_1901 = slice_1900 * slice_1897;
assign slice_6564 = addW_6560[15:0];
assign slice_2657 = mul_2648[17:0];
assign lsl_7320 = mulnw_7319 << 16;
assign slice_3413 = mul_3404[17:0];
assign slice_4169 = addW_4165[17:0];
assign slice_262 = slice_258[17:0];
assign concat_4925 = {concat_4838,slice_4924};
assign add_1018 = lsl_1016 + mul_1017;
assign concat_5681 = {mul_5676,slice_5680};
assign subW_1774 = mul_1773 - mul_1765;
assign slice_6437 = slice_6436[64:32];
assign addW_2530 = concat_2509 + subW_2529;
assign slice_7193 = slice_7192[32:16];
assign mulnw_3286 = slice_3285 * slice_3282;
assign slice_4042 = slice_4033[16:8];
assign slice_135 = mul_134[35:18];
assign slice_4798 = slice_4757[31:0];
assign concat_891 = {addW_889,slice_890};
assign addW_5554 = add_5540 + add_5553;
assign add_1647 = mulnw_1644 + mulnw_1646;
assign add_6310 = mulnw_6307 + mulnw_6309;
assign slice_2403 = addW_2402[33:18];
assign slice_7066 = mul_7065[35:18];
assign subW_3159 = mul_3158 - mul_3150;
assign slice_3915 = slice_3911[15:0];
assign concat_4671 = {mul_4666,slice_4670};
assign mulnw_764 = slice_762 * slice_763;
assign slice_5427 = concat_5381[31:0];
assign subW_1520 = mul_1519 - mul_1511;
assign subW_6183 = subW_6182 - mul_6176;
assign add_2276 = lsl_2274 + mul_2275;
assign add_6939 = lsl_6930 + add_6938;
assign slice_3032 = addW_2990[31:0];
assign add_3788 = lsl_3779 + add_3787;
assign slice_4544 = slice_4534[7:0];
assign concat_637 = {concat_617,slice_636};
assign mulnw_5300 = slice_5299 * slice_5296;
assign subW_1393 = concat_1392 - concat_1220;
assign mulnw_6056 = slice_6055 * slice_6052;
assign concat_2149 = {addW_2147,slice_2148};
assign addW_6812 = concat_6791 + subW_6811;
assign slice_2905 = slice_2904[31:18];
assign mul_7568 = slice_7566 * slice_7567;
assign slice_3661 = slice_3640[31:0];
assign slice_4417 = slice_4416[32:16];
assign mulnw_510 = slice_509 * slice_506;
assign addW_5173 = slice_5168 + slice_5164;
assign slice_1266 = addW_1261[15:0];
assign slice_5929 = slice_5925[17:0];
assign concat_2022 = {addW_2020,slice_2021};
assign slice_6685 = mul_6654[15:0];
assign addW_2778 = slice_2773 + slice_2769;
assign concat_7441 = {mul_7436,slice_7440};
assign lsl_3534 = add_3533 << 8;
assign slice_4290 = slice_4204[63:0];
assign add_383 = lsl_374 + add_382;
assign slice_5046 = concat_4195[255:0];
assign slice_1139 = slice_1138[127:64];
assign add_5802 = mulnw_5799 + mulnw_5801;
assign add_1895 = lsl_1886 + add_1894;
assign addW_6558 = slice_6538 + slice_6519;
assign addW_2651 = slice_2646 + slice_2641;
assign mul_7314 = slice_7312 * slice_7313;
assign addW_3407 = slice_3402 + slice_3398;
assign addW_4163 = slice_4121 + slice_4080;
assign slice_256 = addW_214[31:0];
assign subW_4919 = concat_4918 - concat_4880;
assign mulnw_1012 = slice_1011 * slice_1008;
assign slice_5675 = addW_5674[33:18];
assign mul_1768 = slice_1766 * slice_1767;
assign addW_6431 = slice_6165 + slice_5900;
assign subW_2524 = subW_2523 - mul_2517;
assign concat_7187 = {concat_7100,slice_7186};
assign add_3280 = lsl_3271 + add_3279;
assign mul_4036 = slice_4033 * slice_4035;
assign slice_129 = slice_128[63:32];
assign addW_4792 = add_4778 + add_4791;
assign addW_885 = slice_880 + slice_877;
assign mulnw_5548 = slice_5541 * slice_5547;
assign mulnw_1641 = slice_1639 * slice_1640;
assign mulnw_6304 = slice_6302 * slice_6303;
assign concat_2397 = {addW_2395,slice_2396};
assign slice_7060 = slice_7019[31:0];
assign mul_3153 = slice_3151 * slice_3152;
assign addW_3909 = slice_3643 + slice_3379;
assign slice_4665 = slice_4664[32:16];
assign slice_758 = slice_754[15:0];
assign addW_5421 = concat_5393 + addW_5420;
assign mul_1514 = slice_1512 * slice_1513;
assign slice_6177 = mul_6176[35:18];
assign mulnw_2270 = slice_2269 * slice_2266;
assign slice_6933 = slice_6907[7:0];
assign add_3026 = lsl_3024 + mul_3025;
assign slice_3782 = slice_3772[7:0];
assign slice_4538 = slice_4529[16:8];
assign subW_631 = mul_630 - mul_622;
assign add_5294 = lsl_5285 + add_5293;
assign concat_1387 = {addW_1385,slice_1386};
assign add_6050 = lsl_6041 + add_6049;
assign mul_2143 = slice_2137 * slice_2139;
assign subW_6806 = subW_6805 - mul_6799;
assign subW_2899 = subW_2898 - concat_2855;
assign slice_7562 = addW_7561[33:18];
assign mul_3655 = addW_3653 * addW_3654;
assign add_4411 = lsl_4402 + add_4410;
assign add_504 = lsl_495 + add_503;
assign mul_5167 = slice_5164 * slice_5166;
assign concat_1260 = {concat_1240,slice_1259};
assign slice_5923 = slice_5901[31:0];
assign addW_2016 = slice_2011 + slice_2008;
assign lsl_6679 = add_6678 << 8;
assign mul_2772 = slice_2769 * slice_2771;
assign slice_7435 = slice_7434[31:18];
assign lsl_3528 = mulnw_3527 << 16;
assign addW_4284 = concat_4263 + subW_4283;
assign slice_377 = slice_351[7:0];
assign addW_5040 = concat_4751 + subW_5039;
assign concat_1133 = {addW_1131,slice_1132};
assign mulnw_5796 = slice_5794 * slice_5795;
assign slice_1889 = slice_1879[7:0];
assign subW_6552 = subW_6551 - mul_6545;
assign mul_2645 = slice_2641 * slice_2644;
assign slice_7308 = addW_7307[129:65];
assign mul_3401 = slice_3398 * slice_3400;
assign addW_4157 = add_4143 + add_4156;
assign add_250 = lsl_248 + mul_249;
assign mul_4913 = addW_4911 * addW_4912;
assign concat_1006 = {mul_1001,slice_1005};
assign concat_5669 = {addW_5667,slice_5668};
assign slice_1762 = addW_1761[33:18];
assign subW_6425 = subW_6424 - concat_6336;
assign slice_2518 = mul_2517[35:18];
assign subW_7181 = concat_7180 - concat_7120;
assign slice_3274 = slice_3264[7:0];
assign slice_4030 = concat_4029[63:32];
assign slice_123 = concat_69[31:0];
assign mulnw_4786 = slice_4779 * slice_4785;
assign slice_879 = slice_871[17:0];
assign slice_5542 = slice_5521[16:8];
assign lsl_1635 = add_1634 << 8;
assign slice_6298 = addW_6294[15:0];
assign addW_2391 = slice_2386 + slice_2383;
assign addW_7054 = add_7040 + add_7053;
assign slice_3147 = addW_3146[33:18];
assign slice_3903 = concat_3902[255:128];
assign concat_4659 = {concat_4572,slice_4658};
assign slice_752 = slice_751[32:16];
assign add_5415 = mulnw_5412 + mulnw_5414;
assign slice_1508 = slice_1507[31:18];
assign slice_6171 = slice_6170[63:32];
assign concat_2264 = {mul_2259,slice_2263};
assign slice_6927 = slice_6909[15:8];
assign mulnw_3020 = slice_3019 * slice_3016;
assign slice_3776 = slice_3767[16:8];
assign mul_4532 = slice_4529 * slice_4531;
assign mul_625 = slice_623 * slice_624;
assign slice_5288 = slice_5278[7:0];
assign addW_1381 = slice_1376 + slice_1373;
assign slice_6044 = slice_6034[7:0];
assign slice_2137 = slice_2115[7:0];
assign slice_6800 = mul_6799[35:18];
assign add_2893 = lsl_2884 + add_2892;
assign addW_7556 = concat_7528 + addW_7555;
assign slice_3649 = slice_3645[17:0];
assign slice_4405 = slice_4379[7:0];
assign slice_498 = slice_488[7:0];
assign slice_5161 = mul_5152[17:0];
assign subW_1254 = mul_1253 - mul_1245;
assign mul_5917 = addW_5915 * addW_5916;
assign slice_2010 = slice_2005[17:0];
assign lsl_6673 = mulnw_6672 << 16;
assign slice_2766 = mul_2735[15:0];
assign addW_7429 = concat_7401 + addW_7428;
assign mul_3522 = slice_3516 * slice_3518;
assign subW_4278 = subW_4277 - mul_4271;
assign slice_371 = slice_353[15:8];
assign subW_5034 = subW_5033 - concat_4923;
assign slice_1127 = concat_1103[31:0];
assign slice_5790 = slice_5786[15:0];
assign slice_1883 = slice_1873[16:8];
assign slice_6546 = mul_6545[35:18];
assign slice_2639 = slice_2550[63:0];
assign slice_3395 = mul_3386[17:0];
assign mulnw_4151 = slice_4144 * slice_4150;
assign mulnw_244 = slice_243 * slice_240;
assign slice_4907 = addW_4903[17:0];
assign slice_1000 = addW_999[32:16];
assign addW_5663 = slice_5658 + slice_5655;
assign addW_1756 = concat_1750 + subW_1755;
assign subW_6419 = concat_6418 - concat_6380;
assign addW_2512 = slice_2470 + slice_2430;
assign add_7175 = lsl_7173 + mul_7174;
assign slice_3268 = slice_3258[16:8];
assign mul_4024 = addW_4022 * addW_4023;
assign addW_117 = concat_86 + addW_116;
assign slice_4780 = slice_4759[16:8];
assign slice_873 = slice_27[255:0];
assign add_5536 = mulnw_5533 + mulnw_5535;
assign lsl_1629 = mulnw_1628 << 16;
assign addW_6292 = slice_6272 + slice_6253;
assign slice_2385 = slice_2380[17:0];
assign mulnw_7048 = slice_7041 * slice_7047;
assign addW_3141 = concat_3135 + subW_3140;
assign concat_3897 = {addW_3895,slice_3896};
assign subW_4653 = concat_4652 - concat_4592;
assign slice_746 = concat_745[127:64];
assign mulnw_5409 = slice_5407 * slice_5408;
assign subW_1502 = mul_1501 - mul_1493;
assign slice_6165 = slice_5899[127:0];
assign slice_2258 = slice_2257[32:16];
assign mulnw_6921 = slice_6914 * slice_6920;
assign add_3014 = lsl_3005 + add_3013;
assign mul_3770 = slice_3767 * slice_3769;
assign slice_4526 = concat_4525[63:32];
assign slice_619 = slice_618[31:18];
assign slice_5282 = slice_5273[16:8];
assign slice_1375 = addW_1370[17:0];
assign slice_6038 = slice_6029[16:8];
assign add_2131 = lsl_2129 + mul_2130;
assign addW_6794 = slice_6774 + slice_6734;
assign slice_2887 = slice_2861[7:0];
assign add_7550 = mulnw_7547 + mulnw_7549;
assign slice_3643 = slice_3378[127:0];
assign slice_4399 = slice_4381[15:8];
assign slice_492 = slice_482[16:8];
assign addW_5155 = slice_5150 + slice_5145;
assign mul_1248 = slice_1246 * slice_1247;
assign slice_5911 = slice_5907[17:0];
assign concat_2004 = {addW_2002,slice_2003};
assign mul_6667 = slice_6661 * slice_6663;
assign lsl_2760 = add_2759 << 8;
assign add_7423 = mulnw_7420 + mulnw_7422;
assign slice_3516 = slice_3503[7:0];
assign slice_4272 = mul_4271[35:18];
assign mulnw_365 = slice_358 * slice_364;
assign subW_5028 = concat_5027 - concat_4967;
assign addW_1121 = concat_1115 + subW_1120;
assign slice_5784 = slice_5783[32:16];
assign mul_1877 = slice_1873 * slice_1876;
assign slice_6540 = slice_6521[31:0];
assign concat_2633 = {addW_2631,slice_2632};
assign subW_7296 = subW_7295 - concat_7185;
assign addW_3389 = slice_3384 + slice_3377;
assign slice_4145 = slice_4124[16:8];
assign add_238 = lsl_229 + add_237;
assign addW_4901 = slice_4881 + slice_4840;
assign concat_994 = {addW_992,slice_993};
assign slice_5657 = slice_5652[17:0];
assign concat_1750 = {mul_1745,slice_1749};
assign mul_6413 = addW_6411 * addW_6412;
assign slice_2506 = mul_2475[15:0];
assign mulnw_7169 = slice_7168 * slice_7165;
assign mul_3262 = slice_3258 * slice_3261;
assign slice_4018 = slice_4014[17:0];
assign add_111 = mulnw_108 + mulnw_110;
assign add_4774 = mulnw_4771 + mulnw_4773;
assign concat_867 = {addW_865,slice_866};
assign mulnw_5530 = slice_5528 * slice_5529;
assign mul_1623 = slice_1621 * slice_1622;
assign subW_6286 = subW_6285 - mul_6279;
assign concat_2379 = {addW_2377,slice_2378};
assign slice_7042 = slice_7021[16:8];
assign concat_3135 = {mul_3130,slice_3134};
assign slice_3891 = mul_3882[17:0];
assign add_4647 = lsl_4645 + mul_4646;
assign concat_740 = {addW_738,slice_739};
assign lsl_5403 = add_5402 << 8;
assign mul_1496 = slice_1494 * slice_1495;
assign concat_6159 = {addW_6157,slice_6158};
assign slice_2252 = addW_2251[129:65];
assign slice_6915 = slice_6910[15:8];
assign slice_3008 = slice_2998[7:0];
assign slice_3764 = concat_3763[63:32];
assign mul_4520 = addW_4518 * addW_4519;
assign add_613 = lsl_604 + add_612;
assign mul_5276 = slice_5273 * slice_5275;
assign concat_1369 = {concat_1349,slice_1368};
assign mul_6032 = slice_6029 * slice_6031;
assign mulnw_2125 = slice_2124 * slice_2121;
assign slice_6788 = mul_6779[17:0];
assign slice_2881 = slice_2863[15:8];
assign mulnw_7544 = slice_7542 * slice_7543;
assign slice_3637 = concat_3546[63:0];
assign mulnw_4393 = slice_4386 * slice_4392;
assign mul_486 = slice_482 * slice_485;
assign mul_5149 = slice_5145 * slice_5148;
assign slice_1242 = slice_1241[31:18];
assign slice_5905 = slice_5904[255:128];
assign addW_1998 = slice_1993 + slice_1990;
assign slice_6661 = slice_6648[7:0];
assign lsl_2754 = mulnw_2753 << 16;
assign mulnw_7417 = slice_7415 * slice_7416;
assign slice_3510 = mul_3509[31:16];
assign addW_4266 = slice_4246 + slice_4206;
assign slice_359 = slice_354[15:8];
assign mul_5022 = addW_5020 * addW_5021;
assign concat_1115 = {mul_1110,slice_1114};
assign slice_5778 = concat_5754[31:0];
assign addW_1871 = slice_1784 + slice_1697;
assign subW_6534 = subW_6533 - mul_6527;
assign mul_2627 = slice_2621 * slice_2623;
assign subW_7290 = concat_7289 - concat_7229;
assign mul_3383 = slice_3377 * slice_3382;
assign add_4139 = mulnw_4136 + mulnw_4138;
assign slice_232 = slice_222[7:0];
assign subW_4895 = subW_4894 - mul_4888;
assign addW_988 = slice_983 + slice_980;
assign concat_5651 = {addW_5649,slice_5650};
assign slice_1744 = slice_1743[31:18];
assign slice_6407 = addW_6403[17:0];
assign lsl_2500 = add_2499 << 8;
assign add_7163 = lsl_7154 + add_7162;
assign addW_3256 = slice_3169 + slice_3083;
assign slice_4012 = slice_3992[31:0];
assign mulnw_105 = slice_103 * slice_104;
assign mulnw_4768 = slice_4766 * slice_4767;
assign slice_861 = concat_745[63:0];
assign slice_5524 = slice_5520[15:0];
assign slice_1617 = slice_1616[32:16];
assign slice_6280 = mul_6279[35:18];
assign mul_2373 = slice_2367 * slice_2369;
assign add_7036 = mulnw_7033 + mulnw_7035;
assign slice_3129 = slice_3128[31:18];
assign addW_3885 = slice_3880 + slice_3876;
assign mulnw_4641 = slice_4640 * slice_4637;
assign mul_734 = slice_728 * slice_730;
assign lsl_5397 = mulnw_5396 << 16;
assign slice_1490 = addW_1404[63:0];
assign slice_6153 = mul_6144[17:0];
assign concat_2246 = {addW_2244,slice_2245};
assign slice_6909 = slice_6903[15:0];
assign slice_3002 = slice_2992[16:8];
assign mul_3758 = addW_3756 * addW_3757;
assign slice_4514 = slice_4510[17:0];
assign slice_607 = slice_581[7:0];
assign slice_5270 = mul_5239[15:0];
assign subW_1363 = mul_1362 - mul_1354;
assign slice_6026 = concat_6025[63:32];
assign concat_2119 = {mul_2114,slice_2118};
assign addW_6782 = slice_6777 + slice_6773;
assign mulnw_2875 = slice_2868 * slice_2874;
assign lsl_7538 = add_7537 << 8;
assign addW_3631 = concat_3610 + subW_3630;
assign slice_4387 = slice_4382[15:8];
assign addW_480 = slice_393 + slice_307;
assign slice_5143 = slice_5054[63:0];
assign subW_1236 = mul_1235 - mul_1227;
assign slice_5899 = addW_5052[255:0];
assign slice_1992 = slice_1985[17:0];
assign slice_6655 = mul_6654[31:16];
assign mul_2748 = slice_2742 * slice_2744;
assign lsl_7411 = add_7410 << 8;
assign addW_3504 = slice_3484 + slice_3466;
assign slice_4260 = mul_4251[17:0];
assign slice_353 = addW_348[15:0];
assign slice_5016 = addW_5012[17:0];
assign slice_1109 = addW_1108[33:18];
assign addW_5772 = concat_5766 + subW_5771;
assign subW_1865 = subW_1864 - concat_1821;
assign slice_6528 = mul_6527[35:18];
assign slice_2621 = slice_2599[7:0];
assign mul_7284 = addW_7282 * addW_7283;
assign slice_3377 = slice_3376[31:18];
assign mulnw_4133 = slice_4131 * slice_4132;
assign slice_226 = slice_216[16:8];
assign slice_4889 = mul_4888[35:18];
assign slice_982 = slice_977[17:0];
assign mul_5645 = slice_5639 * slice_5641;
assign addW_1738 = concat_1710 + addW_1737;
assign addW_6401 = slice_6381 + slice_6340;
assign lsl_2494 = mulnw_2493 << 16;
assign slice_7157 = slice_7147[7:0];
assign subW_3250 = subW_3249 - concat_3206;
assign mul_4006 = addW_4004 * addW_4005;
assign lsl_99 = add_98 << 8;
assign slice_4762 = slice_4758[15:0];
assign addW_855 = concat_833 + subW_854;
assign slice_5518 = slice_5517[32:16];
assign add_1611 = lsl_1602 + add_1610;
assign slice_6274 = slice_6255[31:0];
assign slice_2367 = slice_2345[7:0];
assign mulnw_7030 = slice_7028 * slice_7029;
assign addW_3123 = concat_3095 + addW_3122;
assign mul_3879 = slice_3876 * slice_3878;
assign add_4635 = lsl_4626 + add_4634;
assign slice_728 = slice_706[7:0];
assign mul_5391 = slice_5389 * slice_5390;
assign addW_1484 = concat_1463 + subW_1483;
assign addW_6147 = slice_6142 + slice_6138;
assign slice_2240 = concat_2216[31:0];
assign slice_6903 = addW_6902[65:33];
assign mul_2996 = slice_2992 * slice_2995;
assign slice_3752 = slice_3748[17:0];
assign slice_4508 = slice_4487[31:0];
assign slice_601 = slice_583[15:8];
assign lsl_5264 = add_5263 << 8;
assign mul_1357 = slice_1355 * slice_1356;
assign mul_6020 = addW_6018 * addW_6019;
assign slice_2113 = addW_2112[32:16];
assign mul_6776 = slice_6773 * slice_6775;
assign slice_2869 = slice_2864[15:8];
assign lsl_7532 = mulnw_7531 << 16;
assign subW_3625 = subW_3624 - mul_3618;
assign slice_4381 = slice_4375[15:0];
assign subW_474 = subW_473 - concat_430;
assign concat_5137 = {addW_5135,slice_5136};
assign mul_1230 = slice_1228 * slice_1229;
assign concat_5893 = {addW_5891,slice_5892};
assign slice_1986 = slice_1985[31:18];
assign slice_6649 = addW_6608[32:0];
assign slice_2742 = slice_2728[7:0];
assign lsl_7405 = mulnw_7404 << 16;
assign slice_3498 = mul_3489[17:0];
assign addW_4254 = slice_4249 + slice_4245;
assign concat_347 = {concat_327,slice_346};
assign addW_5010 = slice_4968 + slice_4927;
assign concat_1103 = {addW_1101,slice_1102};
assign concat_5766 = {mul_5761,slice_5765};
assign add_1859 = lsl_1850 + add_1858;
assign slice_6522 = slice_6521[63:32];
assign add_2615 = lsl_2613 + mul_2614;
assign slice_7278 = addW_7274[17:0];
assign slice_3371 = concat_3079[127:0];
assign slice_4127 = slice_4123[15:0];
assign mul_220 = slice_216 * slice_219;
assign slice_4883 = slice_4842[31:0];
assign concat_976 = {addW_974,slice_975};
assign slice_5639 = slice_5617[7:0];
assign add_1732 = mulnw_1729 + mulnw_1731;
assign subW_6395 = subW_6394 - mul_6388;
assign mul_2488 = slice_2482 * slice_2484;
assign slice_7151 = slice_7142[16:8];
assign add_3244 = lsl_3235 + add_3243;
assign slice_4000 = slice_3996[17:0];
assign addW_4756 = slice_4490 + slice_4204;
assign subW_849 = subW_848 - mul_842;
assign slice_5512 = concat_5466[31:0];
assign slice_1605 = slice_1579[7:0];
assign subW_6268 = subW_6267 - mul_6261;
assign add_2361 = lsl_2359 + mul_2360;
assign slice_7024 = slice_7020[15:0];
assign add_3117 = mulnw_3114 + mulnw_3116;
assign slice_3873 = concat_3872[63:32];
assign slice_4629 = slice_4619[7:0];
assign add_722 = lsl_720 + mul_721;
assign slice_5385 = addW_5384[32:16];
assign subW_1478 = subW_1477 - mul_1471;
assign mul_6141 = slice_6138 * slice_6140;
assign addW_2234 = concat_2228 + subW_2233;
assign addW_6897 = concat_6854 + subW_6896;
assign addW_2990 = slice_2903 + slice_2817;
assign slice_3746 = slice_3726[31:0];
assign mul_4502 = addW_4500 * addW_4501;
assign mulnw_595 = slice_588 * slice_594;
assign lsl_5258 = mulnw_5257 << 16;
assign slice_1351 = slice_1350[31:18];
assign slice_6014 = slice_6010[17:0];
assign concat_2107 = {addW_2105,slice_2106};
assign slice_6770 = mul_6739[15:0];
assign slice_2863 = addW_2858[15:0];
assign mul_7526 = slice_7524 * slice_7525;
assign slice_3619 = mul_3618[35:18];
assign slice_4375 = addW_4374[65:33];
assign add_468 = lsl_459 + add_467;
assign addW_5131 = slice_5126 + slice_5123;
assign slice_1224 = slice_1138[63:0];
assign slice_5887 = concat_5863[32:0];
assign addW_1980 = concat_1870 + subW_1979;
assign addW_6643 = add_6629 + add_6642;
assign slice_2736 = mul_2735[31:16];
assign mul_7399 = slice_7397 * slice_7398;
assign addW_3492 = slice_3487 + slice_3483;
assign mul_4248 = slice_4245 * slice_4247;
assign subW_341 = mul_340 - mul_332;
assign addW_5004 = add_4990 + add_5003;
assign addW_1097 = slice_1092 + slice_1089;
assign slice_5760 = addW_5759[33:18];
assign slice_1853 = slice_1827[7:0];
assign slice_6516 = concat_6492[31:0];
assign mulnw_2609 = slice_2608 * slice_2605;
assign addW_7272 = slice_7230 + slice_7189;
assign addW_3365 = concat_3255 + subW_3364;
assign slice_4121 = addW_4079[32:0];
assign addW_214 = slice_125 + slice_19;
assign addW_4877 = add_4863 + add_4876;
assign addW_970 = slice_965 + slice_962;
assign add_5633 = lsl_5631 + mul_5632;
assign mulnw_1726 = slice_1724 * slice_1725;
assign slice_6389 = mul_6388[35:18];
assign slice_2482 = slice_2469[7:0];
assign mul_7145 = slice_7142 * slice_7144;
assign slice_3238 = slice_3212[7:0];
assign slice_3994 = slice_3993[31:18];
assign slice_4750 = concat_4749[255:128];
assign slice_843 = mul_842[35:18];
assign addW_5506 = concat_5478 + addW_5505;
assign slice_1599 = slice_1581[15:8];
assign slice_6262 = mul_6261[35:18];
assign mulnw_2355 = slice_2354 * slice_2351;
assign slice_7018 = addW_6731[128:0];
assign mulnw_3111 = slice_3109 * slice_3110;
assign mul_3867 = addW_3865 * addW_3866;
assign slice_4623 = slice_4614[16:8];
assign mulnw_716 = slice_715 * slice_712;
assign addW_5379 = concat_5373 + subW_5378;
assign slice_1472 = mul_1471[35:18];
assign slice_6135 = concat_6134[63:32];
assign concat_2228 = {mul_2223,slice_2227};
assign addW_6891 = add_6877 + add_6890;
assign subW_2984 = subW_2983 - concat_2940;
assign mul_3740 = addW_3738 * addW_3739;
assign slice_4496 = slice_4492[17:0];
assign slice_589 = slice_584[15:8];
assign mul_5252 = slice_5246 * slice_5248;
assign add_1345 = lsl_1336 + add_1344;
assign slice_6008 = slice_5988[31:0];
assign addW_2101 = slice_2096 + slice_2093;
assign lsl_6764 = add_6763 << 8;
assign concat_2857 = {concat_2837,slice_2856};
assign slice_7520 = slice_7519[32:16];
assign addW_3613 = slice_3593 + slice_3553;
assign addW_4369 = concat_4326 + subW_4368;
assign slice_462 = slice_436[7:0];
assign slice_5125 = addW_5120[17:0];
assign addW_1218 = concat_1175 + subW_1217;
assign addW_5881 = concat_5875 + subW_5880;
assign subW_1974 = subW_1973 - concat_1952;
assign mulnw_6637 = slice_6630 * slice_6636;
assign slice_2730 = addW_2729[64:32];
assign slice_7393 = addW_7307[64:0];
assign mul_3486 = slice_3483 * slice_3485;
assign slice_4242 = mul_4211[15:0];
assign mul_335 = slice_333 * slice_334;
assign mulnw_4998 = slice_4991 * slice_4997;
assign slice_1091 = slice_1086[17:0];
assign concat_5754 = {addW_5752,slice_5753};
assign slice_1847 = slice_1829[15:8];
assign addW_6510 = concat_6504 + subW_6509;
assign concat_2603 = {mul_2598,slice_2602};
assign addW_7266 = add_7252 + add_7265;
assign subW_3359 = subW_3358 - concat_3337;
assign add_4115 = lsl_4113 + mul_4114;
assign slice_208 = concat_162[31:0];
assign mulnw_4871 = slice_4864 * slice_4870;
assign slice_964 = slice_958[17:0];
assign mulnw_5627 = slice_5626 * slice_5623;
assign lsl_1720 = add_1719 << 8;
assign slice_6383 = addW_6342[31:0];
assign slice_2476 = mul_2475[31:16];
assign slice_7139 = concat_7138[63:32];
assign slice_3232 = slice_3214[15:8];
assign subW_3988 = subW_3987 - concat_3966;
assign concat_4744 = {addW_4742,slice_4743};
assign addW_837 = slice_794 + slice_754;
assign add_5500 = mulnw_5497 + mulnw_5499;
assign mulnw_1593 = slice_1586 * slice_1592;
assign slice_6256 = slice_6255[63:32];
assign concat_2349 = {mul_2344,slice_2348};
assign slice_7012 = concat_6899[63:0];
assign lsl_3105 = add_3104 << 8;
assign slice_3861 = slice_3857[17:0];
assign mul_4617 = slice_4614 * slice_4616;
assign concat_710 = {mul_705,slice_709};
assign concat_5373 = {mul_5368,slice_5372};
assign addW_1466 = slice_1446 + slice_1406;
assign mul_6129 = addW_6127 * addW_6128;
assign slice_2222 = addW_2221[33:18];
assign mulnw_6885 = slice_6878 * slice_6884;
assign add_2978 = lsl_2969 + add_2977;
assign slice_3734 = slice_3730[17:0];
assign slice_4490 = addW_4203[127:0];
assign slice_583 = slice_576[15:0];
assign slice_5246 = slice_5232[7:0];
assign slice_1339 = slice_1313[7:0];
assign mul_6002 = addW_6000 * addW_6001;
assign slice_2095 = slice_2090[17:0];
assign lsl_6758 = mulnw_6757 << 16;
assign subW_2851 = mul_2850 - mul_2842;
assign add_7514 = lsl_7505 + add_7513;
assign slice_3607 = mul_3598[17:0];
assign addW_4363 = add_4349 + add_4362;
assign slice_456 = slice_438[15:8];
assign concat_5119 = {concat_5099,slice_5118};
assign addW_1212 = add_1198 + add_1211;
assign concat_5875 = {mul_5870,slice_5874};
assign subW_1968 = mul_1967 - mul_1959;
assign slice_6631 = slice_6610[16:8];
assign slice_2724 = concat_2723[127:64];
assign addW_7387 = concat_7366 + subW_7386;
assign slice_3480 = mul_3471[17:0];
assign lsl_4236 = add_4235 << 8;
assign slice_329 = slice_328[31:18];
assign slice_4992 = slice_4971[16:8];
assign concat_1085 = {addW_1083,slice_1084};
assign addW_5748 = slice_5743 + slice_5740;
assign mulnw_1841 = slice_1834 * slice_1840;
assign concat_6504 = {mul_6499,slice_6503};
assign slice_2597 = addW_2596[32:16];
assign mulnw_7260 = slice_7253 * slice_7259;
assign subW_3353 = mul_3352 - mul_3344;
assign mulnw_4109 = slice_4108 * slice_4105;
assign addW_202 = concat_174 + addW_201;
assign slice_4865 = slice_4844[16:8];
assign slice_958 = slice_957[63:32];
assign concat_5621 = {mul_5616,slice_5620};
assign lsl_1714 = mulnw_1713 << 16;
assign addW_6377 = add_6363 + add_6376;
assign slice_2470 = addW_2429[32:0];
assign mul_7133 = addW_7131 * addW_7132;
assign mulnw_3226 = slice_3219 * slice_3225;
assign subW_3982 = mul_3981 - mul_3973;
assign addW_75 = slice_52 + slice_22;
assign slice_4738 = mul_4729[17:0];
assign concat_831 = {addW_829,slice_830};
assign mulnw_5494 = slice_5492 * slice_5493;
assign slice_1587 = slice_1582[15:8];
assign slice_6250 = concat_6204[31:0];
assign slice_2343 = slice_2342[32:16];
assign addW_7006 = concat_6985 + subW_7005;
assign lsl_3099 = mulnw_3098 << 16;
assign slice_3855 = addW_3813[31:0];
assign slice_4611 = concat_4610[63:32];
assign slice_704 = addW_703[32:16];
assign slice_5367 = slice_5366[31:18];
assign slice_1460 = mul_1451[17:0];
assign slice_6123 = slice_6119[17:0];
assign concat_2216 = {addW_2214,slice_2215};
assign slice_6879 = slice_6858[16:8];
assign slice_2972 = slice_2946[7:0];
assign slice_3728 = slice_3727[31:18];
assign slice_4484 = concat_4371[63:0];
assign slice_577 = slice_576[32:16];
assign slice_5240 = mul_5239[31:16];
assign slice_1333 = slice_1315[15:8];
assign slice_5996 = slice_5992[17:0];
assign concat_2089 = {addW_2087,slice_2088};
assign mul_6752 = slice_6746 * slice_6748;
assign mul_2845 = slice_2843 * slice_2844;
assign slice_7508 = slice_7482[7:0];
assign addW_3601 = slice_3596 + slice_3592;
assign mulnw_4357 = slice_4350 * slice_4356;
assign mulnw_450 = slice_443 * slice_449;
assign subW_5113 = mul_5112 - mul_5104;
assign mulnw_1206 = slice_1199 * slice_1205;
assign slice_5869 = addW_5868[33:18];
assign mul_1962 = slice_1960 * slice_1961;
assign add_6625 = mulnw_6622 + mulnw_6624;
assign concat_2718 = {addW_2716,slice_2717};
assign subW_7381 = subW_7380 - mul_7374;
assign addW_3474 = slice_3469 + slice_3464;
assign lsl_4230 = mulnw_4229 << 16;
assign subW_323 = mul_322 - mul_314;
assign add_4986 = mulnw_4983 + mulnw_4985;
assign mul_1079 = slice_1073 * slice_1075;
assign slice_5742 = slice_5737[17:0];
assign slice_1835 = slice_1830[15:8];
assign slice_6498 = addW_6497[33:18];
assign concat_2591 = {addW_2589,slice_2590};
assign slice_7254 = slice_7233[16:8];
assign mul_3347 = slice_3345 * slice_3346;
assign add_4103 = lsl_4094 + add_4102;
assign add_196 = mulnw_193 + mulnw_195;
assign add_4859 = mulnw_4856 + mulnw_4858;
assign subW_952 = concat_951 - concat_891;
assign slice_5615 = slice_5614[32:16];
assign mul_1708 = slice_1706 * slice_1707;
assign mulnw_6371 = slice_6364 * slice_6370;
assign addW_2464 = add_2450 + add_2463;
assign slice_7127 = slice_7123[17:0];
assign slice_3220 = slice_3215[15:8];
assign mul_3976 = slice_3974 * slice_3975;
assign concat_69 = {addW_67,slice_68};
assign addW_4732 = slice_4727 + slice_4723;
assign mul_825 = slice_819 * slice_821;
assign lsl_5488 = add_5487 << 8;
assign slice_1581 = slice_1575[15:0];
assign addW_6244 = concat_6216 + addW_6243;
assign concat_2337 = {addW_2335,slice_2336};
assign subW_7000 = subW_6999 - mul_6993;
assign mul_3093 = slice_3091 * slice_3092;
assign add_3849 = lsl_3847 + mul_3848;
assign mul_4605 = addW_4603 * addW_4604;
assign concat_698 = {addW_696,slice_697};
assign addW_5361 = concat_5355 + subW_5360;
assign addW_1454 = slice_1449 + slice_1445;
assign slice_6117 = addW_6075[31:0];
assign addW_2210 = slice_2205 + slice_2202;
assign add_6873 = mulnw_6870 + mulnw_6872;
assign slice_2966 = slice_2948[15:8];
assign subW_3722 = subW_3721 - concat_3678;
assign addW_4478 = concat_4457 + subW_4477;
assign concat_571 = {concat_305,slice_570};
assign slice_5234 = addW_5233[65:33];
assign mulnw_1327 = slice_1320 * slice_1326;
assign slice_5990 = slice_5989[31:18];
assign addW_2083 = slice_2078 + slice_2075;
assign slice_6746 = slice_6730[7:0];
assign slice_2839 = slice_2838[31:18];
assign slice_7502 = slice_7484[15:8];
assign mul_3595 = slice_3592 * slice_3594;
assign slice_4351 = slice_4330[16:8];
assign slice_444 = slice_439[15:8];
assign mul_5107 = slice_5105 * slice_5106;
assign slice_1200 = slice_1179[16:8];
assign concat_5863 = {addW_5861,slice_5862};
assign slice_1956 = addW_1955[33:18];
assign mulnw_6619 = slice_6617 * slice_6618;
assign mul_2712 = slice_2706 * slice_2708;
assign slice_7375 = mul_7374[35:18];
assign mul_3468 = slice_3464 * slice_3467;
assign mul_4224 = slice_4218 * slice_4220;
assign mul_317 = slice_315 * slice_316;
assign mulnw_4980 = slice_4978 * slice_4979;
assign slice_1073 = slice_1051[7:0];
assign concat_5736 = {addW_5734,slice_5735};
assign slice_1829 = addW_1824[15:0];
assign concat_6492 = {addW_6490,slice_6491};
assign addW_2585 = slice_2580 + slice_2577;
assign add_7248 = mulnw_7245 + mulnw_7247;
assign slice_3341 = addW_3340[33:18];
assign slice_4097 = slice_4087[7:0];
assign mulnw_190 = slice_188 * slice_189;
assign mulnw_4853 = slice_4851 * slice_4852;
assign add_946 = lsl_944 + mul_945;
assign slice_5609 = addW_5608[129:65];
assign slice_1702 = slice_1701[128:64];
assign slice_6365 = slice_6344[16:8];
assign mulnw_2458 = slice_2451 * slice_2457;
assign slice_7121 = slice_7101[31:0];
assign slice_3214 = addW_3209[15:0];
assign slice_3970 = addW_3969[33:18];
assign addW_63 = slice_58 + slice_55;
assign mul_4726 = slice_4723 * slice_4725;
assign slice_819 = slice_797[7:0];
assign lsl_5482 = mulnw_5481 << 16;
assign slice_1575 = addW_1574[65:33];
assign add_6238 = mulnw_6235 + mulnw_6237;
assign slice_2331 = mul_2322[17:0];
assign slice_6994 = mul_6993[35:18];
assign slice_3087 = addW_3086[128:64];
assign mulnw_3843 = slice_3842 * slice_3839;
assign slice_4599 = slice_4595[17:0];
assign addW_692 = slice_687 + slice_684;
assign concat_5355 = {mul_5350,slice_5354};
assign mul_1448 = slice_1445 * slice_1447;
assign add_6111 = lsl_6109 + mul_6110;
assign slice_2204 = slice_2199[17:0];
assign mulnw_6867 = slice_6865 * slice_6866;
assign mulnw_2960 = slice_2953 * slice_2959;
assign add_3716 = lsl_3707 + add_3715;
assign subW_4472 = subW_4471 - mul_4465;
assign subW_565 = concat_564 - concat_392;
assign slice_5228 = concat_5227[127:64];
assign slice_1321 = slice_1316[15:8];
assign subW_5984 = subW_5983 - concat_5940;
assign slice_2077 = slice_2071[17:0];
assign slice_6740 = mul_6739[31:16];
assign subW_2833 = mul_2832 - mul_2824;
assign mulnw_7496 = slice_7489 * slice_7495;
assign slice_3589 = mul_3558[15:0];
assign add_4345 = mulnw_4342 + mulnw_4344;
assign slice_438 = addW_433[15:0];
assign slice_5101 = slice_5100[31:18];
assign add_1194 = mulnw_1191 + mulnw_1193;
assign mul_5857 = slice_5851 * slice_5853;
assign addW_1950 = concat_1922 + addW_1949;
assign slice_6613 = slice_6609[15:0];
assign slice_2706 = slice_2684[7:0];
assign addW_7369 = slice_7349 + slice_7309;
assign slice_3462 = slice_3374[63:0];
assign slice_4218 = slice_4202[7:0];
assign slice_311 = slice_310[127:64];
assign slice_4974 = slice_4970[15:0];
assign add_1067 = lsl_1065 + mul_1066;
assign mul_5730 = slice_5724 * slice_5726;
assign concat_1823 = {concat_1803,slice_1822};
assign addW_6486 = slice_6481 + slice_6478;
assign slice_2579 = slice_2574[17:0];
assign mulnw_7242 = slice_7240 * slice_7241;
assign addW_3335 = concat_3307 + addW_3334;
assign slice_4091 = slice_4081[16:8];
assign lsl_184 = add_183 << 8;
assign slice_4847 = slice_4843[15:0];
assign mulnw_940 = slice_939 * slice_936;
assign addW_5603 = concat_5515 + subW_5602;
assign slice_1696 = addW_1695[256:128];
assign add_6359 = mulnw_6356 + mulnw_6358;
assign slice_2452 = slice_2431[16:8];
assign mul_7115 = addW_7113 * addW_7114;
assign concat_3208 = {concat_3188,slice_3207};
assign addW_3964 = concat_3958 + subW_3963;
assign slice_57 = slice_52[17:0];
assign slice_4720 = concat_4719[63:32];
assign add_813 = lsl_811 + mul_812;
assign mul_5476 = slice_5474 * slice_5475;
assign addW_1569 = concat_1526 + subW_1568;
assign mulnw_6232 = slice_6230 * slice_6231;
assign addW_2325 = slice_2320 + slice_2316;
assign addW_6988 = slice_6946 + slice_6906;
assign concat_3081 = {concat_2815,slice_3080};
assign add_3837 = lsl_3828 + add_3836;
assign slice_4593 = slice_4573[31:0];
assign slice_686 = slice_681[17:0];
assign slice_5349 = slice_5348[31:18];
assign slice_1442 = mul_1411[15:0];
assign mulnw_6105 = slice_6104 * slice_6101;
assign concat_2198 = {addW_2196,slice_2197};
assign slice_6861 = addW_6857[15:0];
assign slice_2954 = slice_2949[15:8];
assign slice_3710 = slice_3684[7:0];
assign slice_4466 = mul_4465[35:18];
assign concat_559 = {addW_557,slice_558};
assign concat_5222 = {addW_5220,slice_5221};
assign slice_1315 = slice_1309[15:0];
assign add_5978 = lsl_5969 + add_5977;
assign slice_2071 = slice_2070[63:32];
assign slice_6734 = slice_6733[64:32];
assign mul_2827 = slice_2825 * slice_2826;
assign slice_7490 = slice_7485[15:8];
assign lsl_3583 = add_3582 << 8;
assign mulnw_4339 = slice_4337 * slice_4338;
assign concat_432 = {concat_412,slice_431};
assign add_5095 = lsl_5086 + add_5094;
assign mulnw_1188 = slice_1186 * slice_1187;
assign slice_5851 = slice_5829[7:0];
assign add_1944 = mulnw_1941 + mulnw_1943;
assign slice_6607 = slice_6606[32:16];
assign add_2700 = lsl_2698 + mul_2699;
assign slice_7363 = mul_7354[17:0];
assign concat_3456 = {addW_3454,slice_3455};
assign slice_4212 = mul_4211[31:16];
assign concat_305 = {addW_303,slice_304};
assign slice_4968 = addW_4926[32:0];
assign mulnw_1061 = slice_1060 * slice_1057;
assign slice_5724 = slice_5702[7:0];
assign subW_1817 = mul_1816 - mul_1808;
assign slice_6480 = slice_6475[17:0];
assign concat_2573 = {addW_2571,slice_2572};
assign slice_7236 = slice_7232[15:0];
assign add_3329 = mulnw_3326 + mulnw_3328;
assign mul_4085 = slice_4081 * slice_4084;
assign lsl_178 = mulnw_177 << 16;
assign slice_4841 = slice_4840[32:16];
assign add_934 = lsl_925 + add_933;
assign subW_5597 = subW_5596 - concat_5575;
assign concat_1690 = {addW_1688,slice_1689};
assign mulnw_6353 = slice_6351 * slice_6352;
assign add_2446 = mulnw_2443 + mulnw_2445;
assign slice_7109 = slice_7105[17:0];
assign subW_3202 = mul_3201 - mul_3193;
assign concat_3958 = {mul_3953,slice_3957};
assign concat_51 = {addW_49,slice_50};
assign mul_4714 = addW_4712 * addW_4713;
assign mulnw_807 = slice_806 * slice_803;
assign slice_5470 = addW_5469[32:16];
assign addW_1563 = add_1549 + add_1562;
assign lsl_6226 = add_6225 << 8;
assign mul_2319 = slice_2316 * slice_2318;
assign slice_6982 = mul_6951[15:0];
assign subW_3075 = concat_3074 - concat_2902;
assign slice_3831 = slice_3821[7:0];
assign mul_4587 = addW_4585 * addW_4586;
assign concat_680 = {addW_678,slice_679};
assign slice_5343 = slice_5342[127:64];
assign lsl_1436 = add_1435 << 8;
assign add_6099 = lsl_6090 + add_6098;
assign mul_2192 = slice_2186 * slice_2188;
assign addW_6855 = slice_6835 + slice_6816;
assign slice_2948 = addW_2943[15:0];
assign slice_3704 = slice_3686[15:8];
assign addW_4460 = slice_4418 + slice_4378;
assign addW_553 = slice_548 + slice_545;
assign mul_5216 = slice_5210 * slice_5212;
assign slice_1309 = addW_1308[64:32];
assign slice_5972 = slice_5946[7:0];
assign subW_2065 = concat_2064 - concat_2004;
assign slice_6728 = slice_6727[128:64];
assign slice_2821 = slice_2820[127:64];
assign slice_7484 = slice_7478[15:0];
assign lsl_3577 = mulnw_3576 << 16;
assign slice_4333 = addW_4329[15:0];
assign subW_426 = mul_425 - mul_417;
assign slice_5089 = slice_5063[7:0];
assign slice_1182 = addW_1178[15:0];
assign add_5845 = lsl_5843 + mul_5844;
assign mulnw_1938 = slice_1936 * slice_1937;
assign slice_6601 = concat_6555[31:0];
assign mulnw_2694 = slice_2693 * slice_2690;
assign addW_7357 = slice_7352 + slice_7348;
assign mul_3450 = slice_3444 * slice_3446;
assign slice_4206 = slice_4205[64:32];
assign slice_299 = concat_273[31:0];
assign add_4962 = lsl_4960 + mul_4961;
assign concat_1055 = {mul_1050,slice_1054};
assign add_5718 = lsl_5716 + mul_5717;
assign mul_1811 = slice_1809 * slice_1810;
assign concat_6474 = {addW_6472,slice_6473};
assign addW_2567 = slice_2562 + slice_2559;
assign slice_7230 = addW_7188[32:0];
assign mulnw_3323 = slice_3321 * slice_3322;
assign addW_4079 = slice_3992 + slice_3906;
assign mul_172 = slice_170 * slice_171;
assign subW_4835 = subW_4834 - concat_4813;
assign slice_928 = slice_918[7:0];
assign subW_5591 = mul_5590 - mul_5582;
assign slice_1684 = concat_1571[63:0];
assign slice_6347 = slice_6343[15:0];
assign mulnw_2440 = slice_2438 * slice_2439;
assign slice_7103 = slice_7102[31:18];
assign mul_3196 = slice_3194 * slice_3195;
assign slice_3952 = slice_3951[31:18];
assign addW_45 = slice_37 + slice_32;
assign slice_4708 = slice_4704[17:0];
assign concat_801 = {mul_796,slice_800};
assign addW_5464 = concat_5458 + subW_5463;
assign mulnw_1557 = slice_1550 * slice_1556;
assign lsl_6220 = mulnw_6219 << 16;
assign slice_2313 = concat_2312[63:32];
assign lsl_6976 = add_6975 << 8;
assign concat_3069 = {addW_3067,slice_3068};
assign slice_3825 = slice_3815[16:8];
assign slice_4581 = slice_4577[17:0];
assign addW_674 = slice_669 + slice_666;
assign subW_5337 = concat_5336 - concat_5142;
assign lsl_1430 = mulnw_1429 << 16;
assign slice_6093 = slice_6083[7:0];
assign slice_2186 = slice_2164[7:0];
assign subW_6849 = subW_6848 - mul_6842;
assign concat_2942 = {concat_2922,slice_2941};
assign mulnw_3698 = slice_3691 * slice_3697;
assign slice_4454 = mul_4423[15:0];
assign slice_547 = addW_542[17:0];
assign slice_5210 = slice_5188[7:0];
assign addW_1303 = concat_1260 + subW_1302;
assign slice_5966 = slice_5948[15:8];
assign add_2059 = lsl_2057 + mul_2058;
assign slice_6722 = concat_6721[511:256];
assign concat_2815 = {addW_2813,slice_2814};
assign slice_7478 = addW_7477[65:33];
assign mul_3571 = slice_3565 * slice_3567;
assign addW_4327 = slice_4307 + slice_4288;
assign mul_420 = slice_418 * slice_419;
assign slice_5083 = slice_5065[15:8];
assign addW_1176 = slice_1156 + slice_1136;
assign mulnw_5839 = slice_5838 * slice_5835;
assign lsl_1932 = add_1931 << 8;
assign addW_6595 = concat_6567 + addW_6594;
assign concat_2688 = {mul_2683,slice_2687};
assign mul_7351 = slice_7348 * slice_7350;
assign slice_3444 = slice_3422[7:0];
assign slice_4200 = slice_4199[128:64];
assign addW_293 = concat_287 + subW_292;
assign mulnw_4956 = slice_4955 * slice_4952;
assign slice_1049 = slice_1048[32:16];
assign mulnw_5712 = slice_5711 * slice_5708;
assign slice_1805 = slice_1804[31:18];
assign mul_6468 = slice_6462 * slice_6464;
assign slice_2561 = slice_2552[17:0];
assign add_7224 = lsl_7222 + mul_7223;
assign lsl_3317 = add_3316 << 8;
assign subW_4073 = subW_4072 - concat_4029;
assign slice_166 = addW_165[32:16];
assign subW_4829 = mul_4828 - mul_4820;
assign slice_922 = slice_913[16:8];
assign mul_5585 = slice_5583 * slice_5584;
assign addW_1678 = concat_1657 + subW_1677;
assign slice_6341 = slice_6340[32:16];
assign slice_2434 = slice_2430[15:0];
assign subW_7097 = subW_7096 - concat_7075;
assign slice_3190 = slice_3189[31:18];
assign addW_3946 = concat_3918 + addW_3945;
assign slice_4702 = addW_4660[31:0];
assign slice_795 = slice_794[32:16];
assign concat_5458 = {mul_5453,slice_5457};
assign slice_1551 = slice_1530[16:8];
assign mul_6214 = slice_6212 * slice_6213;
assign mul_2307 = addW_2305 * addW_2306;
assign lsl_6970 = mulnw_6969 << 16;
assign addW_3063 = slice_3058 + slice_3055;
assign mul_3819 = slice_3815 * slice_3818;
assign slice_4575 = slice_4574[31:18];
assign slice_668 = slice_662[17:0];
assign concat_5331 = {addW_5329,slice_5330};
assign mul_1424 = slice_1418 * slice_1420;
assign slice_6087 = slice_6077[16:8];
assign add_2180 = lsl_2178 + mul_2179;
assign slice_6843 = mul_6842[35:18];
assign subW_2936 = mul_2935 - mul_2927;
assign subW_7599 = concat_7598 - concat_2547;
assign slice_3692 = slice_3687[15:8];
assign lsl_4448 = add_4447 << 8;
assign concat_541 = {concat_521,slice_540};
assign add_5204 = lsl_5202 + mul_5203;
assign addW_1297 = add_1283 + add_1296;
assign mulnw_5960 = slice_5953 * slice_5959;
assign mulnw_2053 = slice_2052 * slice_2049;
assign concat_6716 = {addW_6714,slice_6715};
assign slice_2809 = concat_2785[31:0];
assign addW_7472 = concat_7451 + subW_7471;
assign slice_3565 = slice_3551[7:0];
assign subW_4321 = subW_4320 - mul_4314;
assign slice_414 = slice_413[31:18];
assign mulnw_5077 = slice_5070 * slice_5076;
assign subW_1170 = subW_1169 - mul_1163;
assign concat_5833 = {mul_5828,slice_5832};
assign lsl_1926 = mulnw_1925 << 16;
assign add_6589 = mulnw_6586 + mulnw_6588;
assign slice_2682 = addW_2681[32:16];
assign slice_7345 = mul_7314[15:0];
assign add_3438 = lsl_3436 + mul_3437;
assign slice_4194 = concat_3902[127:0];
assign concat_287 = {mul_282,slice_286};
assign add_4950 = lsl_4941 + add_4949;
assign concat_1043 = {concat_956,slice_1042};
assign concat_5706 = {mul_5701,slice_5705};
assign subW_1799 = mul_1798 - mul_1790;
assign slice_6462 = slice_6440[7:0];
assign slice_2555 = slice_2554[511:256];
assign mulnw_7218 = slice_7217 * slice_7214;
assign lsl_3311 = mulnw_3310 << 16;
assign add_4067 = lsl_4058 + add_4066;
assign addW_160 = concat_154 + subW_159;
assign mul_4823 = slice_4821 * slice_4822;
assign mul_916 = slice_913 * slice_915;
assign slice_5579 = addW_5578[33:18];
assign subW_1672 = subW_1671 - mul_1665;
assign slice_6335 = concat_6289[31:0];
assign slice_2428 = slice_2427[32:16];
assign subW_7091 = mul_7090 - mul_7082;
assign subW_3184 = mul_3183 - mul_3175;
assign add_3940 = mulnw_3937 + mulnw_3939;
assign mul_33 = slice_25 * slice_32;
assign add_4696 = lsl_4694 + mul_4695;
assign addW_789 = concat_761 + addW_788;
assign slice_5452 = slice_5451[31:18];
assign add_1545 = mulnw_1542 + mulnw_1544;
assign slice_6208 = addW_6207[32:16];
assign slice_2301 = slice_2297[17:0];
assign mul_6964 = slice_6958 * slice_6960;
assign slice_3057 = addW_3052[17:0];
assign addW_3813 = slice_3726 + slice_3640;
assign subW_4569 = subW_4568 - concat_4525;
assign slice_662 = slice_661[63:32];
assign addW_5325 = slice_5320 + slice_5317;
assign slice_1418 = slice_1403[7:0];
assign mul_6081 = slice_6077 * slice_6080;
assign mulnw_2174 = slice_2173 * slice_2170;
assign slice_6837 = slice_6818[31:0];
assign mul_2930 = slice_2928 * slice_2929;
assign concat_7593 = {addW_7591,slice_7592};
assign slice_3686 = addW_3681[15:0];
assign lsl_4442 = mulnw_4441 << 16;
assign subW_535 = mul_534 - mul_526;
assign mulnw_5198 = slice_5197 * slice_5194;
assign mulnw_1291 = slice_1284 * slice_1290;
assign slice_5954 = slice_5949[15:8];
assign add_2047 = lsl_2038 + add_2046;
assign slice_6710 = concat_6686[32:0];
assign addW_2803 = concat_2797 + subW_2802;
assign subW_7466 = subW_7465 - mul_7459;
assign slice_3559 = mul_3558[31:16];
assign slice_4315 = mul_4314[35:18];
assign subW_408 = mul_407 - mul_399;
assign slice_5071 = slice_5066[15:8];
assign slice_1164 = mul_1163[35:18];
assign slice_5827 = slice_5826[32:16];
assign mul_1920 = slice_1918 * slice_1919;
assign mulnw_6583 = slice_6581 * slice_6582;
assign concat_2676 = {addW_2674,slice_2675};
assign lsl_7339 = add_7338 << 8;
assign mulnw_3432 = slice_3431 * slice_3428;
assign addW_4188 = concat_4078 + subW_4187;
assign slice_281 = addW_280[33:18];
assign slice_4944 = slice_4934[7:0];
assign subW_1037 = concat_1036 - concat_976;
assign slice_5700 = slice_5699[32:16];
assign mul_1793 = slice_1791 * slice_1792;
assign add_6456 = lsl_6454 + mul_6455;
assign slice_2549 = slice_2548[511:256];
assign add_7212 = lsl_7203 + add_7211;
assign mul_3305 = slice_3303 * slice_3304;
assign slice_4061 = slice_4035[7:0];
assign concat_154 = {mul_149,slice_153};
assign slice_4817 = addW_4816[33:18];
assign slice_910 = concat_909[63:32];
assign addW_5573 = concat_5567 + subW_5572;
assign slice_1666 = mul_1665[35:18];
assign addW_6329 = concat_6301 + addW_6328;
assign concat_2422 = {addW_2420,slice_2421};
assign mul_7085 = slice_7083 * slice_7084;
assign mul_3178 = slice_3176 * slice_3177;
assign mulnw_3934 = slice_3932 * slice_3933;
assign slice_27 = IN2[1023:512];
assign mulnw_4690 = slice_4689 * slice_4686;
assign add_783 = mulnw_780 + mulnw_782;
assign addW_5446 = concat_5440 + subW_5445;
assign mulnw_1539 = slice_1537 * slice_1538;
assign addW_6202 = concat_6196 + subW_6201;
assign slice_2295 = slice_2252[31:0];
assign slice_6958 = slice_6945[7:0];
assign concat_3051 = {concat_3031,slice_3050};
assign subW_3807 = subW_3806 - concat_3763;
assign add_4563 = lsl_4554 + add_4562;
assign subW_656 = concat_655 - concat_617;
assign slice_5319 = addW_5314[17:0];
assign slice_1412 = mul_1411[31:16];
assign addW_6075 = slice_5988 + slice_5901;
assign concat_2168 = {mul_2163,slice_2167};
assign subW_6831 = subW_6830 - mul_6824;
assign slice_2924 = slice_2923[31:18];
assign slice_7587 = concat_7474[64:0];
assign concat_3680 = {concat_3660,slice_3679};
assign mul_4436 = slice_4430 * slice_4432;
assign mul_529 = slice_527 * slice_528;
assign concat_5192 = {mul_5187,slice_5191};
assign slice_1285 = slice_1264[16:8];
assign slice_5948 = addW_5943[15:0];
assign slice_2041 = slice_2031[7:0];
assign addW_6704 = concat_6698 + subW_6703;
assign concat_2797 = {mul_2792,slice_2796};
assign slice_7460 = mul_7459[35:18];
assign slice_3553 = addW_3552[64:32];
assign slice_4309 = slice_4290[31:0];
assign mul_402 = slice_400 * slice_401;
assign slice_5065 = slice_5056[15:0];
assign slice_1158 = slice_1139[31:0];
assign addW_5821 = concat_5793 + addW_5820;
assign slice_1914 = slice_1913[32:16];
assign lsl_6577 = add_6576 << 8;
assign addW_2670 = slice_2665 + slice_2662;
assign lsl_7333 = mulnw_7332 << 16;
assign concat_3426 = {mul_3421,slice_3425};
assign subW_4182 = subW_4181 - concat_4160;
assign concat_275 = {concat_255,slice_274};
assign slice_4938 = slice_4928[16:8];
assign add_1031 = lsl_1029 + mul_1030;
assign concat_5694 = {addW_5692,slice_5693};
assign slice_1787 = slice_1701[63:0];
assign mulnw_6450 = slice_6449 * slice_6446;
assign subW_2543 = concat_2542 - concat_867;
assign slice_7206 = slice_7196[7:0];
assign slice_3299 = slice_3298[32:16];
assign slice_4055 = slice_4037[15:8];
assign slice_148 = slice_147[31:18];
assign addW_4811 = concat_4805 + subW_4810;
assign mul_904 = addW_902 * addW_903;
assign concat_5567 = {mul_5562,slice_5566};
assign addW_1660 = slice_1618 + slice_1578;
assign add_6323 = mulnw_6320 + mulnw_6322;
assign slice_2416 = mul_2407[17:0];
assign slice_7079 = addW_7078[33:18];
assign slice_3172 = addW_3086[63:0];
assign lsl_3928 = add_3927 << 8;
assign add_4684 = lsl_4675 + add_4683;
assign mulnw_777 = slice_775 * slice_776;
assign concat_5440 = {mul_5435,slice_5439};
assign slice_1533 = addW_1529[15:0];
assign concat_6196 = {mul_6191,slice_6195};
assign add_2289 = lsl_2287 + mul_2288;
assign slice_6952 = mul_6951[31:16];
assign subW_3045 = mul_3044 - mul_3036;
assign add_3801 = lsl_3792 + add_3800;
assign slice_4557 = slice_4531[7:0];
assign mul_650 = addW_648 * addW_649;
assign concat_5313 = {concat_5271,slice_5312};
assign slice_1406 = slice_1405[64:32];
assign subW_6069 = subW_6068 - concat_6025;
assign slice_2162 = slice_2161[32:16];
assign slice_6825 = mul_6824[35:18];
assign subW_2918 = mul_2917 - mul_2909;
assign addW_7581 = concat_7560 + subW_7580;
assign subW_3674 = mul_3673 - mul_3665;
assign slice_4430 = slice_4417[7:0];
assign slice_523 = slice_522[31:18];
assign slice_5186 = addW_5185[32:16];
assign add_1279 = mulnw_1276 + mulnw_1278;
assign concat_5942 = {concat_5922,slice_5941};
assign slice_2035 = slice_2026[16:8];
assign concat_6698 = {mul_6693,slice_6697};
assign slice_2791 = addW_2790[33:18];
assign addW_7454 = slice_7434 + slice_7394;
assign slice_3547 = concat_3546[127:64];
assign subW_4303 = subW_4302 - mul_4296;
assign slice_396 = slice_310[63:0];
assign slice_5059 = addW_5058[512:256];
assign subW_1152 = subW_1151 - mul_1145;
assign add_5815 = mulnw_5812 + mulnw_5814;
assign add_1908 = lsl_1899 + add_1907;
assign lsl_6571 = mulnw_6570 << 16;
assign slice_2664 = slice_2659[17:0];
assign mul_7327 = slice_7321 * slice_7323;
assign slice_3420 = addW_3419[32:16];
assign subW_4176 = mul_4175 - mul_4167;
assign subW_269 = mul_268 - mul_260;
assign mul_4932 = slice_4928 * slice_4931;
assign mulnw_1025 = slice_1024 * slice_1021;
assign slice_5688 = mul_5679[17:0];
assign addW_1781 = concat_1760 + subW_1780;
assign concat_6444 = {mul_6439,slice_6443};
assign concat_2537 = {addW_2535,slice_2536};
assign slice_7200 = slice_7190[16:8];
assign add_3293 = lsl_3284 + add_3292;
assign mulnw_4049 = slice_4042 * slice_4048;
assign addW_142 = concat_136 + subW_141;
assign concat_4805 = {mul_4800,slice_4804};
assign slice_898 = slice_894[17:0];
assign slice_5561 = slice_5560[31:18];
assign slice_1654 = mul_1623[15:0];
assign mulnw_6317 = slice_6315 * slice_6316;
assign addW_2410 = slice_2405 + slice_2401;
assign addW_7073 = concat_7067 + subW_7072;
assign addW_3166 = concat_3145 + subW_3165;
assign lsl_3922 = mulnw_3921 << 16;
assign slice_4678 = slice_4668[7:0];
assign lsl_771 = add_770 << 8;
assign slice_5434 = slice_5433[31:18];
assign addW_1527 = slice_1507 + slice_1488;
assign slice_6190 = slice_6189[31:18];
assign mulnw_2283 = slice_2282 * slice_2279;
assign slice_6946 = addW_6905[32:0];
assign mul_3039 = slice_3037 * slice_3038;
assign slice_3795 = slice_3769[7:0];
assign slice_4551 = slice_4533[15:8];
assign slice_644 = addW_640[17:0];
assign add_5307 = lsl_5298 + add_5306;
assign addW_1400 = slice_1134 + slice_869;
assign add_6063 = lsl_6054 + add_6062;
assign concat_2156 = {concat_2069,slice_2155};
assign slice_6819 = slice_6818[63:32];
assign mul_2912 = slice_2910 * slice_2911;
assign subW_7575 = subW_7574 - mul_7568;
assign mul_3668 = slice_3666 * slice_3667;
assign slice_4424 = mul_4423[31:16];
assign add_517 = lsl_508 + add_516;
assign concat_5180 = {addW_5178,slice_5179};
assign mulnw_1273 = slice_1271 * slice_1272;
assign subW_5936 = mul_5935 - mul_5927;
assign mul_2029 = slice_2026 * slice_2028;
assign slice_6692 = addW_6691[33:18];
assign concat_2785 = {addW_2783,slice_2784};
assign slice_7448 = mul_7439[17:0];
assign concat_3541 = {addW_3539,slice_3540};
assign slice_4297 = mul_4296[35:18];
assign addW_390 = concat_347 + subW_389;
assign slice_5053 = addW_5052[512:256];
assign slice_1146 = mul_1145[35:18];
assign mulnw_5809 = slice_5807 * slice_5808;
assign slice_1902 = slice_1876[7:0];
assign mul_6565 = slice_6563 * slice_6564;
assign concat_2658 = {addW_2656,slice_2657};
assign slice_7321 = slice_7306[7:0];
assign concat_3414 = {addW_3412,slice_3413};
assign mul_4170 = slice_4168 * slice_4169;
assign mul_263 = slice_261 * slice_262;
assign addW_4926 = slice_4839 + slice_4753;
assign add_1019 = lsl_1010 + add_1018;
assign addW_5682 = slice_5677 + slice_5673;
assign subW_1775 = subW_1774 - mul_1768;
assign slice_6438 = slice_6437[32:16];
assign slice_2531 = concat_2507[32:0];
assign mul_7194 = slice_7190 * slice_7193;
assign slice_3287 = slice_3261[7:0];
assign slice_4043 = slice_4038[15:8];
assign concat_136 = {mul_131,slice_135};
assign slice_4799 = slice_4798[31:18];
assign slice_892 = slice_870[31:0];
assign addW_5555 = concat_5527 + addW_5554;
assign lsl_1648 = add_1647 << 8;
assign lsl_6311 = add_6310 << 8;
assign mul_2404 = slice_2401 * slice_2403;
assign concat_7067 = {mul_7062,slice_7066};
assign subW_3160 = subW_3159 - mul_3153;
assign mul_3916 = slice_3914 * slice_3915;
assign slice_4672 = slice_4662[16:8];
assign lsl_765 = mulnw_764 << 16;
assign concat_5428 = {addW_5426,slice_5427};
assign subW_1521 = subW_1520 - mul_1514;
assign addW_6184 = concat_6178 + subW_6183;
assign add_2277 = lsl_2268 + add_2276;
assign addW_6940 = add_6926 + add_6939;
assign slice_3033 = slice_3032[31:18];
assign slice_3789 = slice_3771[15:8];
assign mulnw_4545 = slice_4538 * slice_4544;
assign addW_638 = slice_618 + slice_576;
assign slice_5301 = slice_5275[7:0];
assign subW_1394 = subW_1393 - concat_1305;
assign slice_6057 = slice_6031[7:0];
assign subW_2150 = concat_2149 - concat_2089;
assign slice_6813 = concat_6789[31:0];
assign slice_2906 = slice_2820[63:0];
assign slice_7569 = mul_7568[35:18];
assign slice_3662 = slice_3661[31:18];
assign slice_4418 = addW_4377[32:0];
assign slice_511 = slice_485[7:0];
assign addW_5174 = slice_5169 + slice_5166;
assign slice_1267 = addW_1263[15:0];
assign mul_5930 = slice_5928 * slice_5929;
assign slice_2023 = concat_2022[63:32];
assign concat_6686 = {addW_6684,slice_6685};
assign addW_2779 = slice_2774 + slice_2771;
assign addW_7442 = slice_7437 + slice_7433;
assign mul_3535 = slice_3529 * slice_3531;
assign slice_4291 = slice_4290[63:32];
assign addW_384 = add_370 + add_383;
assign concat_5047 = {addW_5045,slice_5046};
assign slice_1140 = slice_1139[63:32];
assign lsl_5803 = add_5802 << 8;
assign slice_1896 = slice_1878[15:8];
assign slice_6559 = addW_6558[32:16];
assign addW_2652 = slice_2647 + slice_2644;
assign slice_7315 = mul_7314[31:16];
assign addW_3408 = slice_3403 + slice_3400;
assign slice_4164 = addW_4163[33:18];
assign slice_257 = slice_256[31:18];
assign subW_4920 = subW_4919 - concat_4898;
assign slice_1013 = slice_1003[7:0];
assign mul_5676 = slice_5673 * slice_5675;
assign slice_1769 = mul_1768[35:18];
assign slice_6432 = addW_6431[128:64];
assign addW_2525 = concat_2519 + subW_2524;
assign addW_7188 = slice_7101 + slice_7015;
assign slice_3281 = slice_3263[15:8];
assign slice_4037 = addW_4032[15:0];
assign slice_130 = slice_129[31:18];
assign addW_4793 = concat_4765 + addW_4792;
assign mul_886 = addW_884 * addW_885;
assign add_5549 = mulnw_5546 + mulnw_5548;
assign lsl_1642 = mulnw_1641 << 16;
assign lsl_6305 = mulnw_6304 << 16;
assign slice_2398 = concat_2397[63:32];
assign slice_7061 = slice_7060[31:18];
assign slice_3154 = mul_3153[35:18];
assign slice_3910 = addW_3909[128:64];
assign mul_4666 = slice_4662 * slice_4665;
assign mul_759 = slice_757 * slice_758;
assign slice_5422 = mul_5391[15:0];
assign slice_1515 = mul_1514[35:18];
assign concat_6178 = {mul_6173,slice_6177};
assign slice_2271 = slice_2261[7:0];
assign mulnw_6934 = slice_6927 * slice_6933;
assign add_3027 = lsl_3018 + add_3026;
assign mulnw_3783 = slice_3776 * slice_3782;
assign slice_4539 = slice_4534[15:8];
assign subW_632 = subW_631 - mul_625;
assign slice_5295 = slice_5277[15:8];
assign subW_1388 = concat_1387 - concat_1349;
assign slice_6051 = slice_6033[15:8];
assign add_2144 = lsl_2142 + mul_2143;
assign addW_6807 = concat_6801 + subW_6806;
assign addW_2900 = concat_2857 + subW_2899;
assign addW_7563 = slice_7521 + slice_7481;
assign subW_3656 = mul_3655 - mul_3647;
assign addW_4412 = add_4398 + add_4411;
assign slice_505 = slice_487[15:8];
assign slice_5168 = slice_5163[17:0];
assign addW_1261 = slice_1241 + slice_1222;
assign slice_5924 = slice_5923[31:18];
assign mul_2017 = addW_2015 * addW_2016;
assign mul_6680 = slice_6674 * slice_6676;
assign slice_2773 = slice_2768[17:0];
assign mul_7436 = slice_7433 * slice_7435;
assign slice_3529 = slice_3507[7:0];
assign slice_4285 = concat_4261[31:0];
assign mulnw_378 = slice_371 * slice_377;
assign slice_5041 = concat_4749[127:0];
assign slice_1134 = slice_868[127:0];
assign lsl_5797 = mulnw_5796 << 16;
assign mulnw_1890 = slice_1883 * slice_1889;
assign addW_6553 = concat_6547 + subW_6552;
assign slice_2646 = slice_2640[17:0];
assign slice_7309 = slice_7308[64:32];
assign slice_3402 = slice_3397[17:0];
assign addW_4158 = concat_4130 + addW_4157;
assign add_251 = lsl_242 + add_250;
assign subW_4914 = mul_4913 - mul_4905;
assign slice_1007 = slice_998[16:8];
assign slice_5670 = concat_5669[63:32];
assign addW_1763 = slice_1743 + slice_1703;
assign addW_6426 = concat_6338 + subW_6425;
assign concat_2519 = {mul_2514,slice_2518};
assign subW_7182 = subW_7181 - concat_7138;
assign mulnw_3275 = slice_3268 * slice_3274;
assign concat_4031 = {concat_4011,slice_4030};
assign concat_124 = {addW_122,slice_123};
assign add_4787 = mulnw_4784 + mulnw_4786;
assign slice_880 = slice_876[17:0];
assign mulnw_5543 = slice_5541 * slice_5542;
assign mul_1636 = slice_1630 * slice_1632;
assign mul_6299 = slice_6297 * slice_6298;
assign mul_2392 = addW_2390 * addW_2391;
assign addW_7055 = concat_7027 + addW_7054;
assign addW_3148 = slice_3128 + slice_3088;
assign concat_3904 = {concat_3638,slice_3903};
assign addW_4660 = slice_4573 + slice_4487;
assign addW_753 = slice_664 + slice_579;
assign lsl_5416 = add_5415 << 8;
assign slice_1509 = slice_1490[31:0];
assign slice_6172 = slice_6171[31:18];
assign slice_2265 = slice_2254[16:8];
assign slice_6928 = slice_6907[16:8];
assign slice_3021 = slice_2995[7:0];
assign slice_3777 = slice_3772[15:8];
assign slice_4533 = addW_4528[15:0];
assign slice_626 = mul_625[35:18];
assign mulnw_5289 = slice_5282 * slice_5288;
assign mul_1382 = addW_1380 * addW_1381;
assign mulnw_6045 = slice_6038 * slice_6044;
assign mulnw_2138 = slice_2137 * slice_2134;
assign concat_6801 = {mul_6796,slice_6800};
assign addW_2894 = add_2880 + add_2893;
assign slice_7557 = mul_7526[15:0];
assign mul_3650 = slice_3648 * slice_3649;
assign mulnw_4406 = slice_4399 * slice_4405;
assign mulnw_499 = slice_492 * slice_498;
assign concat_5162 = {addW_5160,slice_5161};
assign subW_1255 = subW_1254 - mul_1248;
assign subW_5918 = mul_5917 - mul_5909;
assign slice_2011 = slice_2007[17:0];
assign slice_6674 = slice_6652[7:0];
assign concat_2767 = {addW_2765,slice_2766};
assign slice_7430 = mul_7399[15:0];
assign add_3523 = lsl_3521 + mul_3522;
assign addW_4279 = concat_4273 + subW_4278;
assign slice_372 = slice_351[16:8];
assign addW_5035 = concat_4925 + subW_5034;
assign concat_1128 = {addW_1126,slice_1127};
assign mul_5791 = slice_5789 * slice_5790;
assign slice_1884 = slice_1879[15:8];
assign concat_6547 = {mul_6542,slice_6546};
assign slice_2640 = slice_2639[63:32];
assign addW_7303 = slice_7014 + slice_6727;
assign concat_3396 = {addW_3394,slice_3395};
assign add_4152 = mulnw_4149 + mulnw_4151;
assign slice_245 = slice_219[7:0];
assign mul_4908 = slice_4906 * slice_4907;
assign mul_1001 = slice_998 * slice_1000;
assign mul_5664 = addW_5662 * addW_5663;
assign slice_1757 = mul_1748[17:0];
assign subW_6420 = subW_6419 - concat_6398;
assign slice_2513 = addW_2512[33:18];
assign add_7176 = lsl_7167 + add_7175;
assign slice_3269 = slice_3264[15:8];
assign subW_4025 = mul_4024 - mul_4016;
assign slice_118 = mul_84[15:0];
assign mulnw_4781 = slice_4779 * slice_4780;
assign slice_874 = slice_873[255:128];
assign lsl_5537 = add_5536 << 8;
assign slice_1630 = slice_1617[7:0];
assign slice_6293 = addW_6292[32:16];
assign slice_2386 = slice_2382[17:0];
assign add_7049 = mulnw_7046 + mulnw_7048;
assign slice_3142 = mul_3133[17:0];
assign subW_3898 = concat_3897 - concat_3725;
assign subW_4654 = subW_4653 - concat_4610;
assign concat_747 = {concat_660,slice_746};
assign lsl_5410 = mulnw_5409 << 16;
assign subW_1503 = subW_1502 - mul_1496;
assign slice_6166 = slice_6165[127:64];
assign mul_2259 = slice_2254 * slice_2258;
assign add_6922 = mulnw_6919 + mulnw_6921;
assign slice_3015 = slice_2997[15:8];
assign slice_3771 = addW_3766[15:0];
assign concat_4527 = {concat_4507,slice_4526};
assign slice_620 = slice_579[31:0];
assign slice_5283 = slice_5278[15:8];
assign slice_1376 = addW_1372[17:0];
assign slice_6039 = slice_6034[15:8];
assign add_2132 = lsl_2123 + add_2131;
assign slice_6795 = addW_6794[33:18];
assign mulnw_2888 = slice_2881 * slice_2887;
assign lsl_7551 = add_7550 << 8;
assign slice_3644 = slice_3643[127:64];
assign slice_4400 = slice_4379[16:8];
assign slice_493 = slice_488[15:8];
assign addW_5156 = slice_5151 + slice_5148;
assign slice_1249 = mul_1248[35:18];
assign mul_5912 = slice_5910 * slice_5911;
assign slice_2005 = slice_1984[31:0];
assign add_6668 = lsl_6666 + mul_6667;
assign mul_2761 = slice_2755 * slice_2757;
assign lsl_7424 = add_7423 << 8;
assign mulnw_3517 = slice_3516 * slice_3513;
assign concat_4273 = {mul_4268,slice_4272};
assign add_366 = mulnw_363 + mulnw_365;
assign subW_5029 = subW_5028 - concat_5007;
assign slice_1122 = mul_1113[17:0];
assign addW_5785 = slice_5698 + slice_5613;
assign slice_1878 = slice_1872[15:0];
assign slice_6541 = slice_6540[31:18];
assign subW_2634 = concat_2633 - concat_2573;
assign addW_7297 = concat_7187 + subW_7296;
assign addW_3390 = slice_3385 + slice_3382;
assign mulnw_4146 = slice_4144 * slice_4145;
assign slice_239 = slice_221[15:8];
assign slice_4902 = addW_4901[33:18];
assign slice_995 = concat_994[63:32];
assign slice_5658 = slice_5654[17:0];
assign addW_1751 = slice_1746 + slice_1742;
assign subW_6414 = mul_6413 - mul_6405;
assign concat_2507 = {addW_2505,slice_2506};
assign slice_7170 = slice_7144[7:0];
assign slice_3263 = slice_3257[15:0];
assign mul_4019 = slice_4017 * slice_4018;
assign lsl_112 = add_111 << 8;
assign lsl_4775 = add_4774 << 8;
assign slice_868 = slice_10[255:0];
assign lsl_5531 = mulnw_5530 << 16;
assign slice_1624 = mul_1623[31:16];
assign addW_6287 = concat_6281 + subW_6286;
assign slice_2380 = slice_2338[31:0];
assign mulnw_7043 = slice_7041 * slice_7042;
assign addW_3136 = slice_3131 + slice_3127;
assign concat_3892 = {addW_3890,slice_3891};
assign add_4648 = lsl_4639 + add_4647;
assign subW_741 = concat_740 - concat_680;
assign mul_5404 = slice_5398 * slice_5400;
assign slice_1497 = mul_1496[35:18];
assign subW_6160 = concat_6159 - concat_5987;
assign slice_2253 = slice_2252[64:32];
assign mulnw_6916 = slice_6914 * slice_6915;
assign mulnw_3009 = slice_3002 * slice_3008;
assign concat_3765 = {concat_3745,slice_3764};
assign subW_4521 = mul_4520 - mul_4512;
assign addW_614 = add_600 + add_613;
assign slice_5277 = slice_5272[15:0];
assign addW_1370 = slice_1350 + slice_1309;
assign slice_6033 = addW_6028[15:0];
assign slice_2126 = slice_2116[7:0];
assign concat_6789 = {addW_6787,slice_6788};
assign slice_2882 = slice_2861[16:8];
assign lsl_7545 = mulnw_7544 << 16;
assign concat_3638 = {addW_3636,slice_3637};
assign add_4394 = mulnw_4391 + mulnw_4393;
assign slice_487 = slice_481[15:0];
assign slice_5150 = slice_5144[17:0];
assign slice_1243 = slice_1224[31:0];
assign slice_5906 = slice_5905[127:64];
assign mul_1999 = addW_1997 * addW_1998;
assign mulnw_6662 = slice_6661 * slice_6658;
assign slice_2755 = slice_2733[7:0];
assign lsl_7418 = mulnw_7417 << 16;
assign concat_3511 = {mul_3506,slice_3510};
assign slice_4267 = addW_4266[33:18];
assign mulnw_360 = slice_358 * slice_359;
assign subW_5023 = mul_5022 - mul_5014;
assign addW_1116 = slice_1111 + slice_1107;
assign concat_5779 = {addW_5777,slice_5778};
assign slice_1872 = addW_1871[65:33];
assign addW_6535 = concat_6529 + subW_6534;
assign add_2628 = lsl_2626 + mul_2627;
assign subW_7291 = subW_7290 - concat_7269;
assign slice_3384 = slice_3376[17:0];
assign lsl_4140 = add_4139 << 8;
assign mulnw_233 = slice_226 * slice_232;
assign addW_4896 = concat_4890 + subW_4895;
assign mul_989 = addW_987 * addW_988;
assign slice_5652 = slice_5609[31:0];
assign mul_1745 = slice_1742 * slice_1744;
assign mul_6408 = slice_6406 * slice_6407;
assign mul_2501 = slice_2495 * slice_2497;
assign slice_7164 = slice_7146[15:8];
assign slice_3257 = addW_3256[65:33];
assign slice_4013 = slice_4012[31:18];
assign lsl_106 = mulnw_105 << 16;
assign lsl_4769 = mulnw_4768 << 16;
assign concat_862 = {addW_860,slice_861};
assign mul_5525 = slice_5523 * slice_5524;
assign slice_1618 = addW_1577[32:0];
assign concat_6281 = {mul_6276,slice_6280};
assign add_2374 = lsl_2372 + mul_2373;
assign lsl_7037 = add_7036 << 8;
assign mul_3130 = slice_3127 * slice_3129;
assign addW_3886 = slice_3881 + slice_3878;
assign slice_4642 = slice_4616[7:0];
assign add_735 = lsl_733 + mul_734;
assign slice_5398 = slice_5385[7:0];
assign slice_1491 = slice_1490[63:32];
assign concat_6154 = {addW_6152,slice_6153};
assign slice_2247 = concat_2246[255:128];
assign slice_6910 = slice_6906[15:0];
assign slice_3003 = slice_2998[15:8];
assign subW_3759 = mul_3758 - mul_3750;
assign mul_4515 = slice_4513 * slice_4514;
assign mulnw_608 = slice_601 * slice_607;
assign concat_5271 = {addW_5269,slice_5270};
assign subW_1364 = subW_1363 - mul_1357;
assign concat_6027 = {concat_6007,slice_6026};
assign slice_2120 = slice_2111[16:8];
assign addW_6783 = slice_6778 + slice_6775;
assign add_2876 = mulnw_2873 + mulnw_2875;
assign mul_7539 = slice_7533 * slice_7535;
assign slice_3632 = concat_3608[31:0];
assign mulnw_4388 = slice_4386 * slice_4387;
assign slice_481 = addW_480[64:32];
assign slice_5144 = slice_5143[63:32];
assign subW_1237 = subW_1236 - mul_1230;
assign slice_5900 = slice_5899[255:128];
assign slice_1993 = slice_1989[17:0];
assign concat_6656 = {mul_6651,slice_6655};
assign add_2749 = lsl_2747 + mul_2748;
assign mul_7412 = slice_7406 * slice_7408;
assign slice_3505 = addW_3504[32:16];
assign concat_4261 = {addW_4259,slice_4260};
assign slice_354 = addW_350[15:0];
assign mul_5017 = slice_5015 * slice_5016;
assign mul_1110 = slice_1107 * slice_1109;
assign slice_5773 = mul_5764[17:0];
assign addW_1866 = concat_1823 + subW_1865;
assign concat_6529 = {mul_6524,slice_6528};
assign mulnw_2622 = slice_2621 * slice_2618;
assign subW_7285 = mul_7284 - mul_7276;
assign slice_3378 = slice_2554[255:0];
assign lsl_4134 = mulnw_4133 << 16;
assign slice_227 = slice_222[15:8];
assign concat_4890 = {mul_4885,slice_4889};
assign slice_983 = slice_979[17:0];
assign add_5646 = lsl_5644 + mul_5645;
assign slice_1739 = mul_1708[15:0];
assign slice_6402 = addW_6401[33:18];
assign slice_2495 = slice_2473[7:0];
assign mulnw_7158 = slice_7151 * slice_7157;
assign addW_3251 = concat_3208 + subW_3250;
assign subW_4007 = mul_4006 - mul_3998;
assign mul_100 = slice_94 * slice_96;
assign mul_4763 = slice_4761 * slice_4762;
assign slice_856 = concat_831[32:0];
assign addW_5519 = slice_5432 + slice_5347;
assign addW_1612 = add_1598 + add_1611;
assign slice_6275 = slice_6274[31:18];
assign mulnw_2368 = slice_2367 * slice_2364;
assign lsl_7031 = mulnw_7030 << 16;
assign slice_3124 = mul_3093[15:0];
assign slice_3880 = addW_3875[17:0];
assign slice_4636 = slice_4618[15:8];
assign mulnw_729 = slice_728 * slice_725;
assign slice_5392 = mul_5391[31:16];
assign slice_1485 = concat_1461[31:0];
assign addW_6148 = slice_6143 + slice_6140;
assign concat_2241 = {addW_2239,slice_2240};
assign slice_6904 = slice_6903[32:16];
assign slice_2997 = slice_2991[15:0];
assign mul_3753 = slice_3751 * slice_3752;
assign slice_4509 = slice_4508[31:18];
assign slice_602 = slice_581[16:8];
assign mul_5265 = slice_5259 * slice_5261;
assign slice_1358 = mul_1357[35:18];
assign subW_6021 = mul_6020 - mul_6012;
assign mul_2114 = slice_2111 * slice_2113;
assign slice_6777 = slice_6772[17:0];
assign mulnw_2870 = slice_2868 * slice_2869;
assign slice_7533 = slice_7520[7:0];
assign addW_3626 = concat_3620 + subW_3625;
assign slice_4382 = slice_4378[15:0];
assign addW_475 = concat_432 + subW_474;
assign subW_5138 = concat_5137 - concat_5099;
assign slice_1231 = mul_1230[35:18];
assign subW_5894 = concat_5893 - concat_5341;
assign slice_1987 = addW_1700[127:0];
assign slice_6650 = slice_6649[32:16];
assign mulnw_2743 = slice_2742 * slice_2739;
assign slice_7406 = slice_7392[7:0];
assign concat_3499 = {addW_3497,slice_3498};
assign addW_4255 = slice_4250 + slice_4247;
assign addW_348 = slice_328 + slice_308;
assign slice_5011 = addW_5010[33:18];
assign slice_1104 = concat_1103[63:32];
assign addW_5767 = slice_5762 + slice_5758;
assign addW_1860 = add_1846 + add_1859;
assign slice_6523 = slice_6522[31:18];
assign add_2616 = lsl_2607 + add_2615;
assign mul_7279 = slice_7277 * slice_7278;
assign concat_3372 = {addW_3370,slice_3371};
assign mul_4128 = slice_4126 * slice_4127;
assign slice_221 = slice_215[15:0];
assign slice_4884 = slice_4883[31:18];
assign slice_977 = slice_957[31:0];
assign mulnw_5640 = slice_5639 * slice_5636;
assign lsl_1733 = add_1732 << 8;
assign addW_6396 = concat_6390 + subW_6395;
assign add_2489 = lsl_2487 + mul_2488;
assign slice_7152 = slice_7147[15:8];
assign addW_3245 = add_3231 + add_3244;
assign mul_4001 = slice_3999 * slice_4000;
assign slice_94 = slice_77[7:0];
assign slice_4757 = addW_4756[129:65];
assign addW_850 = concat_844 + subW_849;
assign concat_5513 = {addW_5511,slice_5512};
assign mulnw_1606 = slice_1599 * slice_1605;
assign addW_6269 = concat_6263 + subW_6268;
assign add_2362 = lsl_2353 + add_2361;
assign mul_7025 = slice_7023 * slice_7024;
assign lsl_3118 = add_3117 << 8;
assign concat_3874 = {concat_3854,slice_3873};
assign mulnw_4630 = slice_4623 * slice_4629;
assign add_723 = lsl_714 + add_722;
assign addW_5386 = slice_5366 + slice_5348;
assign addW_1479 = concat_1473 + subW_1478;
assign slice_6142 = addW_6137[17:0];
assign slice_2235 = mul_2226[17:0];
assign slice_6898 = concat_6852[31:0];
assign slice_2991 = addW_2990[64:32];
assign slice_3747 = slice_3746[31:18];
assign subW_4503 = mul_4502 - mul_4494;
assign add_596 = mulnw_593 + mulnw_595;
assign slice_5259 = slice_5237[7:0];
assign slice_1352 = addW_1311[31:0];
assign mul_6015 = slice_6013 * slice_6014;
assign slice_2108 = concat_2107[63:32];
assign concat_6771 = {addW_6769,slice_6770};
assign slice_2864 = addW_2860[15:0];
assign slice_7527 = mul_7526[31:16];
assign concat_3620 = {mul_3615,slice_3619};
assign slice_4376 = slice_4375[32:16];
assign addW_469 = add_455 + add_468;
assign mul_5132 = addW_5130 * addW_5131;
assign slice_1225 = slice_1224[63:32];
assign concat_5888 = {addW_5886,slice_5887};
assign slice_1981 = concat_1868[63:0];
assign addW_6644 = concat_6616 + addW_6643;
assign concat_2737 = {mul_2732,slice_2736};
assign slice_7400 = mul_7399[31:16];
assign addW_3493 = slice_3488 + slice_3485;
assign slice_4249 = slice_4244[17:0];
assign subW_342 = subW_341 - mul_335;
assign addW_5005 = concat_4977 + addW_5004;
assign mul_1098 = addW_1096 * addW_1097;
assign mul_5761 = slice_5758 * slice_5760;
assign mulnw_1854 = slice_1847 * slice_1853;
assign concat_6517 = {addW_6515,slice_6516};
assign slice_2610 = slice_2600[7:0];
assign slice_7273 = addW_7272[33:18];
assign slice_3366 = concat_3253[63:0];
assign slice_4122 = slice_4121[32:16];
assign slice_215 = addW_214[64:32];
assign addW_4878 = concat_4850 + addW_4877;
assign mul_971 = addW_969 * addW_970;
assign add_5634 = lsl_5625 + add_5633;
assign lsl_1727 = mulnw_1726 << 16;
assign concat_6390 = {mul_6385,slice_6389};
assign mulnw_2483 = slice_2482 * slice_2479;
assign slice_7146 = addW_7141[15:0];
assign mulnw_3239 = slice_3232 * slice_3238;
assign slice_3995 = addW_3909[63:0];
assign concat_4751 = {concat_4485,slice_4750};
assign concat_844 = {mul_839,slice_843};
assign slice_5507 = mul_5476[15:0];
assign slice_1600 = slice_1579[16:8];
assign concat_6263 = {mul_6258,slice_6262};
assign slice_2356 = slice_2346[7:0];
assign slice_7019 = slice_7018[128:64];
assign lsl_3112 = mulnw_3111 << 16;
assign subW_3868 = mul_3867 - mul_3859;
assign slice_4624 = slice_4619[15:8];
assign slice_717 = slice_707[7:0];
assign slice_5380 = mul_5371[17:0];
assign concat_1473 = {mul_1468,slice_1472};
assign concat_6136 = {concat_6116,slice_6135};
assign addW_2229 = slice_2224 + slice_2220;
assign addW_6892 = concat_6864 + addW_6891;
assign addW_2985 = concat_2942 + subW_2984;
assign subW_3741 = mul_3740 - mul_3732;
assign mul_4497 = slice_4495 * slice_4496;
assign mulnw_590 = slice_588 * slice_589;
assign add_5253 = lsl_5251 + mul_5252;
assign addW_1346 = add_1332 + add_1345;
assign slice_6009 = slice_6008[31:18];
assign mul_2102 = addW_2100 * addW_2101;
assign mul_6765 = slice_6759 * slice_6761;
assign addW_2858 = slice_2838 + slice_2818;
assign slice_7521 = addW_7480[32:0];
assign slice_3614 = addW_3613[33:18];
assign slice_4370 = concat_4324[31:0];
assign mulnw_463 = slice_456 * slice_462;
assign slice_5126 = addW_5122[17:0];
assign slice_1219 = concat_1173[31:0];
assign slice_5882 = mul_5873[17:0];
assign addW_1975 = concat_1954 + subW_1974;
assign add_6638 = mulnw_6635 + mulnw_6637;
assign slice_2731 = slice_2730[32:16];
assign slice_7394 = slice_7393[64:32];
assign slice_3487 = slice_3482[17:0];
assign concat_4243 = {addW_4241,slice_4242};
assign slice_336 = mul_335[35:18];
assign add_4999 = mulnw_4996 + mulnw_4998;
assign slice_1092 = slice_1088[17:0];
assign slice_5755 = concat_5754[63:32];
assign slice_1848 = slice_1827[16:8];
assign slice_6511 = mul_6502[17:0];
assign slice_2604 = slice_2595[16:8];
assign addW_7267 = concat_7239 + addW_7266;
assign addW_3360 = concat_3339 + subW_3359;
assign add_4116 = lsl_4107 + add_4115;
assign concat_209 = {addW_207,slice_208};
assign add_4872 = mulnw_4869 + mulnw_4871;
assign slice_965 = slice_961[17:0];
assign slice_5628 = slice_5618[7:0];
assign mul_1721 = slice_1715 * slice_1717;
assign slice_6384 = slice_6383[31:18];
assign concat_2477 = {mul_2472,slice_2476};
assign concat_7140 = {concat_7120,slice_7139};
assign slice_3233 = slice_3212[16:8];
assign addW_3989 = concat_3968 + subW_3988;
assign slice_82 = addW_75[15:0];
assign subW_4745 = concat_4744 - concat_4572;
assign slice_838 = addW_837[33:18];
assign lsl_5501 = add_5500 << 8;
assign add_1594 = mulnw_1591 + mulnw_1593;
assign slice_6257 = slice_6256[31:18];
assign slice_2350 = slice_2340[16:8];
assign concat_7013 = {addW_7011,slice_7012};
assign mul_3106 = slice_3100 * slice_3102;
assign mul_3862 = slice_3860 * slice_3861;
assign slice_4618 = addW_4613[15:0];
assign slice_711 = slice_702[16:8];
assign addW_5374 = slice_5369 + slice_5365;
assign slice_1467 = addW_1466[33:18];
assign subW_6130 = mul_6129 - mul_6121;
assign mul_2223 = slice_2220 * slice_2222;
assign add_6886 = mulnw_6883 + mulnw_6885;
assign addW_2979 = add_2965 + add_2978;
assign mul_3735 = slice_3733 * slice_3734;
assign slice_4491 = slice_4490[127:64];
assign slice_584 = slice_580[15:0];
assign mulnw_5247 = slice_5246 * slice_5243;
assign mulnw_1340 = slice_1333 * slice_1339;
assign subW_6003 = mul_6002 - mul_5994;
assign slice_2096 = slice_2092[17:0];
assign slice_6759 = slice_6737[7:0];
assign subW_2852 = subW_2851 - mul_2845;
assign addW_7515 = add_7501 + add_7514;
assign concat_3608 = {addW_3606,slice_3607};
assign addW_4364 = concat_4336 + addW_4363;
assign slice_457 = slice_436[16:8];
assign addW_5120 = slice_5100 + slice_5056;
assign addW_1213 = concat_1185 + addW_1212;
assign addW_5876 = slice_5871 + slice_5867;
assign subW_1969 = subW_1968 - mul_1962;
assign mulnw_6632 = slice_6630 * slice_6631;
assign concat_2725 = {concat_2638,slice_2724};
assign slice_7388 = concat_7364[31:0];
assign concat_3481 = {addW_3479,slice_3480};
assign mul_4237 = slice_4231 * slice_4233;
assign slice_330 = slice_311[31:0];
assign mulnw_4993 = slice_4991 * slice_4992;
assign slice_1086 = addW_1044[31:0];
assign mul_5749 = addW_5747 * addW_5748;
assign add_1842 = mulnw_1839 + mulnw_1841;
assign addW_6505 = slice_6500 + slice_6496;
assign mul_2598 = slice_2595 * slice_2597;
assign add_7261 = mulnw_7258 + mulnw_7260;
assign subW_3354 = subW_3353 - mul_3347;
assign slice_4110 = slice_4084[7:0];
assign slice_203 = mul_172[15:0];
assign mulnw_4866 = slice_4864 * slice_4865;
assign slice_959 = slice_958[31:18];
assign slice_5622 = slice_5611[16:8];
assign slice_1715 = slice_1699[7:0];
assign addW_6378 = concat_6350 + addW_6377;
assign slice_2471 = slice_2470[32:16];
assign subW_7134 = mul_7133 - mul_7125;
assign add_3227 = mulnw_3224 + mulnw_3226;
assign subW_3983 = subW_3982 - mul_3976;
assign concat_4739 = {addW_4737,slice_4738};
assign slice_832 = concat_831[65:33];
assign lsl_5495 = mulnw_5494 << 16;
assign mulnw_1588 = slice_1586 * slice_1587;
assign concat_6251 = {addW_6249,slice_6250};
assign mul_2344 = slice_2340 * slice_2343;
assign slice_7007 = concat_6983[32:0];
assign slice_3100 = slice_3085[7:0];
assign slice_3856 = slice_3855[31:18];
assign concat_4612 = {concat_4592,slice_4611};
assign mul_705 = slice_702 * slice_704;
assign mul_5368 = slice_5365 * slice_5367;
assign concat_1461 = {addW_1459,slice_1460};
assign mul_6124 = slice_6122 * slice_6123;
assign slice_2217 = concat_2216[63:32];
assign mulnw_6880 = slice_6878 * slice_6879;
assign mulnw_2973 = slice_2966 * slice_2972;
assign slice_3729 = slice_3643[63:0];
assign concat_4485 = {addW_4483,slice_4484};
assign addW_578 = slice_310 + slice_29;
assign concat_5241 = {mul_5236,slice_5240};
assign slice_1334 = slice_1313[16:8];
assign mul_5997 = slice_5995 * slice_5996;
assign slice_2090 = slice_2070[31:0];
assign add_6753 = lsl_6751 + mul_6752;
assign slice_2846 = mul_2845[35:18];
assign mulnw_7509 = slice_7502 * slice_7508;
assign addW_3602 = slice_3597 + slice_3594;
assign add_4358 = mulnw_4355 + mulnw_4357;
assign add_451 = mulnw_448 + mulnw_450;
assign subW_5114 = subW_5113 - mul_5107;
assign add_1207 = mulnw_1204 + mulnw_1206;
assign mul_5870 = slice_5867 * slice_5869;
assign slice_1963 = mul_1962[35:18];
assign lsl_6626 = add_6625 << 8;
assign subW_2719 = concat_2718 - concat_2658;
assign addW_7382 = concat_7376 + subW_7381;
assign addW_3475 = slice_3470 + slice_3467;
assign slice_4231 = slice_4209[7:0];
assign subW_324 = subW_323 - mul_317;
assign lsl_4987 = add_4986 << 8;
assign add_1080 = lsl_1078 + mul_1079;
assign slice_5743 = slice_5739[17:0];
assign mulnw_1836 = slice_1834 * slice_1835;
assign mul_6499 = slice_6496 * slice_6498;
assign slice_2592 = concat_2591[63:32];
assign mulnw_7255 = slice_7253 * slice_7254;
assign slice_3348 = mul_3347[35:18];
assign slice_4104 = slice_4086[15:8];
assign lsl_197 = add_196 << 8;
assign lsl_4860 = add_4859 << 8;
assign subW_953 = subW_952 - concat_909;
assign mul_5616 = slice_5611 * slice_5615;
assign slice_1709 = mul_1708[31:16];
assign add_6372 = mulnw_6369 + mulnw_6371;
assign addW_2465 = concat_2437 + addW_2464;
assign mul_7128 = slice_7126 * slice_7127;
assign mulnw_3221 = slice_3219 * slice_3220;
assign slice_3977 = mul_3976[35:18];
assign slice_70 = concat_69[63:32];
assign addW_4733 = slice_4728 + slice_4725;
assign add_826 = lsl_824 + mul_825;
assign mul_5489 = slice_5483 * slice_5485;
assign slice_1582 = slice_1578[15:0];
assign slice_6245 = mul_6214[15:0];
assign slice_2338 = addW_2251[64:0];
assign addW_7001 = concat_6995 + subW_7000;
assign slice_3094 = mul_3093[31:16];
assign add_3850 = lsl_3841 + add_3849;
assign subW_4606 = mul_4605 - mul_4597;
assign slice_699 = concat_698[63:32];
assign slice_5362 = mul_5353[17:0];
assign addW_1455 = slice_1450 + slice_1447;
assign slice_6118 = slice_6117[31:18];
assign mul_2211 = addW_2209 * addW_2210;
assign lsl_6874 = add_6873 << 8;
assign slice_2967 = slice_2946[16:8];
assign addW_3723 = concat_3680 + subW_3722;
assign slice_4479 = concat_4455[32:0];
assign slice_5235 = slice_5234[32:16];
assign add_1328 = mulnw_1325 + mulnw_1327;
assign slice_5991 = slice_5905[63:0];
assign mul_2084 = addW_2082 * addW_2083;
assign mulnw_6747 = slice_6746 * slice_6743;
assign slice_2840 = slice_2821[31:0];
assign slice_7503 = slice_7482[16:8];
assign slice_3596 = slice_3591[17:0];
assign mulnw_4352 = slice_4350 * slice_4351;
assign mulnw_445 = slice_443 * slice_444;
assign slice_5108 = mul_5107[35:18];
assign mulnw_1201 = slice_1199 * slice_1200;
assign slice_5864 = concat_5863[65:33];
assign addW_1957 = slice_1915 + slice_1875;
assign lsl_6620 = mulnw_6619 << 16;
assign add_2713 = lsl_2711 + mul_2712;
assign concat_7376 = {mul_7371,slice_7375};
assign slice_3469 = slice_3463[17:0];
assign add_4225 = lsl_4223 + mul_4224;
assign slice_318 = mul_317[35:18];
assign lsl_4981 = mulnw_4980 << 16;
assign mulnw_1074 = slice_1073 * slice_1070;
assign slice_5737 = slice_5695[31:0];
assign slice_1830 = addW_1826[15:0];
assign slice_6493 = concat_6492[63:32];
assign mul_2586 = addW_2584 * addW_2585;
assign lsl_7249 = add_7248 << 8;
assign addW_3342 = slice_3300 + slice_3260;
assign mulnw_4098 = slice_4091 * slice_4097;
assign lsl_191 = mulnw_190 << 16;
assign lsl_4854 = mulnw_4853 << 16;
assign add_947 = lsl_938 + add_946;
assign slice_5610 = slice_5609[64:32];
assign slice_1703 = slice_1702[64:32];
assign mulnw_6366 = slice_6364 * slice_6365;
assign add_2459 = mulnw_2456 + mulnw_2458;
assign slice_7122 = slice_7121[31:18];
assign slice_3215 = addW_3211[15:0];
assign addW_3971 = slice_3951 + slice_3911;
assign mul_64 = addW_62 * addW_63;
assign slice_4727 = addW_4722[17:0];
assign mulnw_820 = slice_819 * slice_816;
assign slice_5483 = slice_5470[7:0];
assign slice_1576 = slice_1575[32:16];
assign lsl_6239 = add_6238 << 8;
assign concat_2332 = {addW_2330,slice_2331};
assign concat_6995 = {mul_6990,slice_6994};
assign slice_3088 = slice_3087[64:32];
assign slice_3844 = slice_3818[7:0];
assign mul_4600 = slice_4598 * slice_4599;
assign mul_693 = addW_691 * addW_692;
assign addW_5356 = slice_5351 + slice_5345;
assign slice_1449 = slice_1444[17:0];
assign add_6112 = lsl_6103 + add_6111;
assign slice_2205 = slice_2201[17:0];
assign lsl_6868 = mulnw_6867 << 16;
assign add_2961 = mulnw_2958 + mulnw_2960;
assign addW_3717 = add_3703 + add_3716;
assign addW_4473 = concat_4467 + subW_4472;
assign subW_566 = subW_565 - concat_477;
assign concat_5229 = {concat_5142,slice_5228};
assign mulnw_1322 = slice_1320 * slice_1321;
assign addW_5985 = concat_5942 + subW_5984;
assign slice_2078 = slice_2074[17:0];
assign concat_6741 = {mul_6736,slice_6740};
assign subW_2834 = subW_2833 - mul_2827;
assign add_7497 = mulnw_7494 + mulnw_7496;
assign concat_3590 = {addW_3588,slice_3589};
assign lsl_4346 = add_4345 << 8;
assign slice_439 = addW_435[15:0];
assign slice_5102 = slice_5061[31:0];
assign lsl_1195 = add_1194 << 8;
assign add_5858 = lsl_5856 + mul_5857;
assign slice_1951 = mul_1920[15:0];
assign mul_6614 = slice_6612 * slice_6613;
assign mulnw_2707 = slice_2706 * slice_2703;
assign slice_7370 = addW_7369[33:18];
assign slice_3463 = slice_3462[63:32];
assign mulnw_4219 = slice_4218 * slice_4215;
assign slice_312 = slice_311[63:32];
assign mul_4975 = slice_4973 * slice_4974;
assign add_1068 = lsl_1059 + add_1067;
assign add_5731 = lsl_5729 + mul_5730;
assign addW_1824 = slice_1804 + slice_1785;
assign mul_6487 = addW_6485 * addW_6486;
assign slice_2580 = slice_2576[17:0];
assign lsl_7243 = mulnw_7242 << 16;
assign slice_3336 = mul_3305[15:0];
assign slice_4092 = slice_4087[15:8];
assign mul_185 = slice_179 * slice_181;
assign mul_4848 = slice_4846 * slice_4847;
assign slice_941 = slice_915[7:0];
assign slice_5604 = concat_5513[63:0];
assign slice_1697 = slice_1696[128:64];
assign lsl_6360 = add_6359 << 8;
assign mulnw_2453 = slice_2451 * slice_2452;
assign subW_7116 = mul_7115 - mul_7107;
assign addW_3209 = slice_3189 + slice_3170;
assign slice_3965 = mul_3956[17:0];
assign slice_58 = slice_54[17:0];
assign concat_4721 = {concat_4701,slice_4720};
assign add_814 = lsl_805 + add_813;
assign slice_5477 = mul_5476[31:16];
assign slice_1570 = concat_1524[31:0];
assign lsl_6233 = mulnw_6232 << 16;
assign addW_2326 = slice_2321 + slice_2318;
assign slice_6989 = addW_6988[33:18];
assign addW_3082 = slice_2816 + slice_2550;
assign slice_3838 = slice_3820[15:8];
assign slice_4594 = slice_4593[31:18];
assign slice_687 = slice_683[17:0];
assign mul_5350 = slice_5345 * slice_5349;
assign concat_1443 = {addW_1441,slice_1442};
assign slice_6106 = slice_6080[7:0];
assign slice_2199 = addW_2157[31:0];
assign mul_6862 = slice_6860 * slice_6861;
assign mulnw_2955 = slice_2953 * slice_2954;
assign mulnw_3711 = slice_3704 * slice_3710;
assign concat_4467 = {mul_4462,slice_4466};
assign subW_560 = concat_559 - concat_521;
assign subW_5223 = concat_5222 - concat_5162;
assign slice_1316 = slice_1312[15:0];
assign addW_5979 = add_5965 + add_5978;
assign slice_2072 = slice_2071[31:18];
assign slice_6735 = slice_6734[32:16];
assign slice_2828 = mul_2827[35:18];
assign mulnw_7491 = slice_7489 * slice_7490;
assign mul_3584 = slice_3578 * slice_3580;
assign lsl_4340 = mulnw_4339 << 16;
assign addW_433 = slice_413 + slice_394;
assign addW_5096 = add_5082 + add_5095;
assign lsl_1189 = mulnw_1188 << 16;
assign mulnw_5852 = slice_5851 * slice_5848;
assign lsl_1945 = add_1944 << 8;
assign addW_6608 = slice_6521 + slice_6436;
assign add_2701 = lsl_2692 + add_2700;
assign concat_7364 = {addW_7362,slice_7363};
assign subW_3457 = concat_3456 - concat_3396;
assign concat_4213 = {mul_4208,slice_4212};
assign slice_306 = slice_13[127:0];
assign slice_4969 = slice_4968[32:16];
assign slice_1062 = slice_1052[7:0];
assign mulnw_5725 = slice_5724 * slice_5721;
assign subW_1818 = subW_1817 - mul_1811;
assign slice_6481 = slice_6477[17:0];
assign slice_2574 = slice_2551[31:0];
assign mul_7237 = slice_7235 * slice_7236;
assign lsl_3330 = add_3329 << 8;
assign slice_4086 = slice_4080[15:0];
assign slice_179 = slice_166[7:0];
assign slice_4842 = addW_4756[64:0];
assign slice_935 = slice_917[15:8];
assign addW_5598 = concat_5577 + subW_5597;
assign slice_1691 = concat_1690[511:256];
assign lsl_6354 = mulnw_6353 << 16;
assign lsl_2447 = add_2446 << 8;
assign mul_7110 = slice_7108 * slice_7109;
assign subW_3203 = subW_3202 - mul_3196;
assign addW_3959 = slice_3954 + slice_3950;
assign slice_52 = slice_19[31:0];
assign subW_4715 = mul_4714 - mul_4706;
assign slice_808 = slice_798[7:0];
assign addW_5471 = slice_5451 + slice_5433;
assign addW_1564 = concat_1536 + addW_1563;
assign mul_6227 = slice_6221 * slice_6223;
assign slice_2320 = addW_2315[17:0];
assign concat_6983 = {addW_6981,slice_6982};
assign subW_3076 = subW_3075 - concat_2987;
assign mulnw_3832 = slice_3825 * slice_3831;
assign subW_4588 = mul_4587 - mul_4579;
assign slice_681 = slice_661[31:0];
assign slice_5344 = slice_5343[63:32];
assign mul_1437 = slice_1431 * slice_1433;
assign slice_6100 = slice_6082[15:8];
assign add_2193 = lsl_2191 + mul_2192;
assign slice_6856 = addW_6855[32:16];
assign slice_2949 = addW_2945[15:0];
assign slice_3705 = slice_3684[16:8];
assign slice_4461 = addW_4460[33:18];
assign mul_554 = addW_552 * addW_553;
assign add_5217 = lsl_5215 + mul_5216;
assign slice_1310 = slice_1309[32:16];
assign mulnw_5973 = slice_5966 * slice_5972;
assign subW_2066 = subW_2065 - concat_2022;
assign slice_6729 = slice_6728[64:32];
assign slice_2822 = slice_2821[63:32];
assign slice_7485 = slice_7481[15:0];
assign slice_3578 = slice_3556[7:0];
assign mul_4334 = slice_4332 * slice_4333;
assign subW_427 = subW_426 - mul_420;
assign mulnw_5090 = slice_5083 * slice_5089;
assign mul_1183 = slice_1181 * slice_1182;
assign add_5846 = lsl_5837 + add_5845;
assign lsl_1939 = mulnw_1938 << 16;
assign concat_6602 = {addW_6600,slice_6601};
assign slice_2695 = slice_2685[7:0];
assign addW_7358 = slice_7353 + slice_7350;
assign add_3451 = lsl_3449 + mul_3450;
assign slice_4207 = slice_4206[32:16];
assign concat_300 = {addW_298,slice_299};
assign add_4963 = lsl_4954 + add_4962;
assign slice_1056 = slice_1046[16:8];
assign add_5719 = lsl_5710 + add_5718;
assign slice_1812 = mul_1811[35:18];
assign slice_6475 = slice_6432[31:0];
assign mul_2568 = addW_2566 * addW_2567;
assign slice_7231 = slice_7230[32:16];
assign lsl_3324 = mulnw_3323 << 16;
assign slice_4080 = addW_4079[65:33];
assign slice_173 = mul_172[31:16];
assign addW_4836 = concat_4815 + subW_4835;
assign mulnw_929 = slice_922 * slice_928;
assign subW_5592 = subW_5591 - mul_5585;
assign concat_1685 = {addW_1683,slice_1684};
assign mul_6348 = slice_6346 * slice_6347;
assign lsl_2441 = mulnw_2440 << 16;
assign slice_7104 = slice_7018[63:0];
assign slice_3197 = mul_3196[35:18];
assign mul_3953 = slice_3950 * slice_3952;
assign mul_46 = addW_44 * addW_45;
assign mul_4709 = slice_4707 * slice_4708;
assign slice_802 = slice_793[16:8];
assign slice_5465 = mul_5456[17:0];
assign add_1558 = mulnw_1555 + mulnw_1557;
assign slice_6221 = slice_6208[7:0];
assign concat_2314 = {concat_2294,slice_2313};
assign mul_6977 = slice_6971 * slice_6973;
assign subW_3070 = concat_3069 - concat_3031;
assign slice_3826 = slice_3821[15:8];
assign mul_4582 = slice_4580 * slice_4581;
assign mul_675 = addW_673 * addW_674;
assign subW_5338 = subW_5337 - concat_5227;
assign slice_1431 = slice_1409[7:0];
assign mulnw_6094 = slice_6087 * slice_6093;
assign mulnw_2187 = slice_2186 * slice_2183;
assign addW_6850 = concat_6844 + subW_6849;
assign addW_2943 = slice_2923 + slice_2904;
assign add_3699 = mulnw_3696 + mulnw_3698;
assign concat_4455 = {addW_4453,slice_4454};
assign slice_548 = addW_544[17:0];
assign mulnw_5211 = slice_5210 * slice_5207;
assign slice_1304 = concat_1258[31:0];
assign slice_5967 = slice_5946[16:8];
assign add_2060 = lsl_2051 + add_2059;
assign concat_6723 = {concat_5898,slice_6722};
assign slice_2816 = slice_2549[127:0];
assign slice_7479 = slice_7478[32:16];
assign add_3572 = lsl_3570 + mul_3571;
assign slice_4328 = addW_4327[32:16];
assign slice_421 = mul_420[35:18];
assign slice_5084 = slice_5063[16:8];
assign slice_1177 = addW_1176[32:16];
assign slice_5840 = slice_5830[7:0];
assign mul_1933 = slice_1927 * slice_1929;
assign slice_6596 = mul_6565[15:0];
assign slice_2689 = slice_2680[16:8];
assign slice_7352 = slice_7347[17:0];
assign mulnw_3445 = slice_3444 * slice_3441;
assign slice_4201 = slice_4200[64:32];
assign slice_294 = mul_285[17:0];
assign slice_4957 = slice_4931[7:0];
assign mul_1050 = slice_1046 * slice_1049;
assign slice_5713 = slice_5703[7:0];
assign slice_1806 = slice_1787[31:0];
assign add_6469 = lsl_6467 + mul_6468;
assign slice_2562 = slice_2558[17:0];
assign add_7225 = lsl_7216 + add_7224;
assign mul_3318 = slice_3312 * slice_3314;
assign addW_4074 = concat_4031 + subW_4073;
assign addW_167 = slice_147 + slice_129;
assign subW_4830 = subW_4829 - mul_4823;
assign slice_923 = slice_918[15:8];
assign slice_5586 = mul_5585[35:18];
assign slice_1679 = concat_1655[32:0];
assign addW_6342 = slice_6255 + slice_6170;
assign mul_2435 = slice_2433 * slice_2434;
assign addW_7098 = concat_7077 + subW_7097;
assign slice_3191 = slice_3172[31:0];
assign slice_3947 = mul_3916[15:0];
assign slice_40 = mul_38[35:18];
assign slice_4703 = slice_4702[31:18];
assign mul_796 = slice_793 * slice_795;
assign addW_5459 = slice_5454 + slice_5450;
assign mulnw_1552 = slice_1550 * slice_1551;
assign slice_6215 = mul_6214[31:16];
assign subW_2308 = mul_2307 - mul_2299;
assign slice_6971 = slice_6949[7:0];
assign mul_3064 = addW_3062 * addW_3063;
assign slice_3820 = slice_3814[15:0];
assign slice_4576 = slice_4490[63:0];
assign slice_669 = slice_665[17:0];
assign subW_5332 = concat_5331 - concat_5271;
assign add_1425 = lsl_1423 + mul_1424;
assign slice_6088 = slice_6083[15:8];
assign add_2181 = lsl_2172 + add_2180;
assign concat_6844 = {mul_6839,slice_6843};
assign subW_2937 = subW_2936 - mul_2930;
assign subW_7600 = subW_7599 - concat_5047;
assign mulnw_3693 = slice_3691 * slice_3692;
assign mul_4449 = slice_4443 * slice_4445;
assign addW_542 = slice_522 + slice_481;
assign add_5205 = lsl_5196 + add_5204;
assign addW_1298 = concat_1270 + addW_1297;
assign add_5961 = mulnw_5958 + mulnw_5960;
assign slice_2054 = slice_2028[7:0];
assign subW_6717 = concat_6716 - concat_6164;
assign concat_2810 = {addW_2808,slice_2809};
assign slice_7473 = concat_7449[31:0];
assign mulnw_3566 = slice_3565 * slice_3562;
assign addW_4322 = concat_4316 + subW_4321;
assign slice_415 = slice_396[31:0];
assign add_5078 = mulnw_5075 + mulnw_5077;
assign addW_1171 = concat_1165 + subW_1170;
assign slice_5834 = slice_5825[16:8];
assign slice_1927 = slice_1914[7:0];
assign lsl_6590 = add_6589 << 8;
assign mul_2683 = slice_2680 * slice_2682;
assign concat_7346 = {addW_7344,slice_7345};
assign add_3439 = lsl_3430 + add_3438;
assign concat_4195 = {addW_4193,slice_4194};
assign addW_288 = slice_283 + slice_279;
assign slice_4951 = slice_4933[15:8];
assign addW_1044 = slice_957 + slice_870;
assign slice_5707 = slice_5697[16:8];
assign subW_1800 = subW_1799 - mul_1793;
assign mulnw_6463 = slice_6462 * slice_6459;
assign slice_2556 = slice_2555[255:128];
assign slice_7219 = slice_7193[7:0];
assign slice_3312 = slice_3299[7:0];
assign addW_4068 = add_4054 + add_4067;
assign slice_161 = mul_152[17:0];
assign slice_4824 = mul_4823[35:18];
assign slice_917 = addW_912[15:0];
assign addW_5580 = slice_5560 + slice_5520;
assign addW_1673 = concat_1667 + subW_1672;
assign concat_6336 = {addW_6334,slice_6335};
assign addW_2429 = slice_2341 + slice_2256;
assign subW_7092 = subW_7091 - mul_7085;
assign subW_3185 = subW_3184 - mul_3178;
assign lsl_3941 = add_3940 << 8;
assign add_4697 = lsl_4688 + add_4696;
assign slice_790 = mul_759[15:0];
assign mul_5453 = slice_5450 * slice_5452;
assign lsl_1546 = add_1545 << 8;
assign addW_6209 = slice_6189 + slice_6171;
assign mul_2302 = slice_2300 * slice_2301;
assign add_6965 = lsl_6963 + mul_6964;
assign slice_3058 = addW_3054[17:0];
assign slice_3814 = addW_3813[64:32];
assign addW_4570 = concat_4527 + subW_4569;
assign slice_663 = slice_662[31:18];
assign mul_5326 = addW_5324 * addW_5325;
assign mulnw_1419 = slice_1418 * slice_1415;
assign slice_6082 = slice_6076[15:0];
assign slice_2175 = slice_2165[7:0];
assign slice_6838 = slice_6837[31:18];
assign slice_2931 = mul_2930[35:18];
assign subW_7594 = concat_7593 - concat_5898;
assign slice_3687 = addW_3683[15:0];
assign slice_4443 = slice_4421[7:0];
assign subW_536 = subW_535 - mul_529;
assign slice_5199 = slice_5189[7:0];
assign add_1292 = mulnw_1289 + mulnw_1291;
assign mulnw_5955 = slice_5953 * slice_5954;
assign slice_2048 = slice_2030[15:8];
assign concat_6711 = {addW_6709,slice_6710};
assign slice_2804 = mul_2795[17:0];
assign addW_7467 = concat_7461 + subW_7466;
assign concat_3560 = {mul_3555,slice_3559};
assign concat_4316 = {mul_4311,slice_4315};
assign subW_409 = subW_408 - mul_402;
assign mulnw_5072 = slice_5070 * slice_5071;
assign concat_1165 = {mul_1160,slice_1164};
assign mul_5828 = slice_5825 * slice_5827;
assign slice_1921 = mul_1920[31:16];
assign lsl_6584 = mulnw_6583 << 16;
assign slice_2677 = concat_2676[63:32];
assign mul_7340 = slice_7334 * slice_7336;
assign slice_3433 = slice_3423[7:0];
assign slice_4189 = concat_4076[63:0];
assign mul_282 = slice_279 * slice_281;
assign mulnw_4945 = slice_4938 * slice_4944;
assign subW_1038 = subW_1037 - concat_994;
assign mul_5701 = slice_5697 * slice_5700;
assign slice_1794 = mul_1793[35:18];
assign add_6457 = lsl_6448 + add_6456;
assign slice_2550 = slice_2549[255:128];
assign slice_7213 = slice_7195[15:8];
assign slice_3306 = mul_3305[31:16];
assign mulnw_4062 = slice_4055 * slice_4061;
assign addW_155 = slice_150 + slice_146;
assign addW_4818 = slice_4798 + slice_4758;
assign concat_911 = {concat_891,slice_910};
assign slice_5574 = mul_5565[17:0];
assign concat_1667 = {mul_1662,slice_1666};
assign slice_6330 = mul_6299[15:0];
assign slice_2423 = concat_2422[129:65];
assign slice_7086 = mul_7085[35:18];
assign slice_3179 = mul_3178[35:18];
assign lsl_3935 = mulnw_3934 << 16;
assign slice_28 = slice_27[511:256];
assign slice_4691 = slice_4665[7:0];
assign lsl_784 = add_783 << 8;
assign slice_5447 = mul_5438[17:0];
assign lsl_1540 = mulnw_1539 << 16;
assign slice_6203 = mul_6194[17:0];
assign slice_2296 = slice_2295[31:18];
assign mulnw_6959 = slice_6958 * slice_6955;
assign addW_3052 = slice_3032 + slice_2991;
assign addW_3808 = concat_3765 + subW_3807;
assign addW_4564 = add_4550 + add_4563;
assign subW_657 = subW_656 - concat_635;
assign slice_5320 = addW_5316[17:0];
assign concat_1413 = {mul_1408,slice_1412};
assign slice_6076 = addW_6075[64:32];
assign slice_2169 = slice_2159[16:8];
assign addW_6832 = concat_6826 + subW_6831;
assign slice_2925 = slice_2906[31:0];
assign concat_7588 = {addW_7586,slice_7587};
assign addW_3681 = slice_3661 + slice_3641;
assign add_4437 = lsl_4435 + mul_4436;
assign slice_530 = mul_529[35:18];
assign slice_5193 = slice_5184[16:8];
assign mulnw_1286 = slice_1284 * slice_1285;
assign slice_5949 = addW_5945[15:0];
assign mulnw_2042 = slice_2035 * slice_2041;
assign slice_6705 = mul_6696[17:0];
assign addW_2798 = slice_2793 + slice_2789;
assign concat_7461 = {mul_7456,slice_7460};
assign slice_3554 = slice_3553[32:16];
assign slice_4310 = slice_4309[31:18];
assign slice_403 = mul_402[35:18];
assign slice_5066 = slice_5062[15:0];
assign slice_1159 = slice_1158[31:18];
assign slice_5822 = mul_5791[15:0];
assign slice_1915 = addW_1874[32:0];
assign mul_6578 = slice_6572 * slice_6574;
assign mul_2671 = addW_2669 * addW_2670;
assign slice_7334 = slice_7312[7:0];
assign slice_3427 = slice_3418[16:8];
assign addW_4183 = concat_4162 + subW_4182;
assign slice_4939 = slice_4934[15:8];
assign add_1032 = lsl_1023 + add_1031;
assign slice_5695 = addW_5608[64:0];
assign slice_1788 = slice_1787[63:32];
assign slice_6451 = slice_6441[7:0];
assign subW_2544 = subW_2543 - concat_1690;
assign mulnw_7207 = slice_7200 * slice_7206;
assign slice_3300 = addW_3259[32:0];
assign slice_4056 = slice_4035[16:8];
assign mul_149 = slice_146 * slice_148;
assign slice_4812 = mul_4803[17:0];
assign subW_905 = mul_904 - mul_896;
assign addW_5568 = slice_5563 + slice_5559;
assign slice_1661 = addW_1660[33:18];
assign lsl_6324 = add_6323 << 8;
assign concat_2417 = {addW_2415,slice_2416};
assign addW_7080 = slice_7060 + slice_7020;
assign slice_3173 = slice_3172[63:32];
assign mul_3929 = slice_3923 * slice_3925;
assign slice_22 = slice_19[63:32];
assign slice_4685 = slice_4667[15:8];
assign lsl_778 = mulnw_777 << 16;
assign addW_5441 = slice_5436 + slice_5431;
assign mul_1534 = slice_1532 * slice_1533;
assign addW_6197 = slice_6192 + slice_6188;
assign add_2290 = lsl_2281 + add_2289;
assign concat_6953 = {mul_6948,slice_6952};
assign subW_3046 = subW_3045 - mul_3039;
assign addW_3802 = add_3788 + add_3801;
assign mulnw_4558 = slice_4551 * slice_4557;
assign subW_651 = mul_650 - mul_642;
assign addW_5314 = slice_5272 + slice_5231;
assign slice_1407 = slice_1406[32:16];
assign addW_6070 = concat_6027 + subW_6069;
assign mul_2163 = slice_2159 * slice_2162;
assign concat_6826 = {mul_6821,slice_6825};
assign subW_2919 = subW_2918 - mul_2912;
assign slice_7582 = concat_7558[32:0];
assign subW_3675 = subW_3674 - mul_3668;
assign mulnw_4431 = slice_4430 * slice_4427;
assign slice_524 = addW_483[31:0];
assign mul_5187 = slice_5184 * slice_5186;
assign lsl_1280 = add_1279 << 8;
assign addW_5943 = slice_5923 + slice_5902;
assign slice_2036 = slice_2031[15:8];
assign addW_6699 = slice_6694 + slice_6690;
assign mul_2792 = slice_2789 * slice_2791;
assign slice_7455 = addW_7454[33:18];
assign concat_3548 = {concat_3461,slice_3547};
assign addW_4304 = concat_4298 + subW_4303;
assign slice_397 = slice_396[63:32];
assign slice_5060 = slice_5059[256:128];
assign addW_1153 = concat_1147 + subW_1152;
assign lsl_5816 = add_5815 << 8;
assign addW_1909 = add_1895 + add_1908;
assign slice_6572 = slice_6559[7:0];
assign slice_2665 = slice_2661[17:0];
assign add_7328 = lsl_7326 + mul_7327;
assign mul_3421 = slice_3418 * slice_3420;
assign subW_4177 = subW_4176 - mul_4170;
assign subW_270 = subW_269 - mul_263;
assign slice_4933 = slice_4927[15:0];
assign slice_1026 = slice_1000[7:0];
assign concat_5689 = {addW_5687,slice_5688};
assign slice_1782 = concat_1758[31:0];
assign slice_6445 = slice_6434[16:8];
assign subW_2538 = concat_2537 - concat_1982;
assign slice_7201 = slice_7196[15:8];
assign addW_3294 = add_3280 + add_3293;
assign add_4050 = mulnw_4047 + mulnw_4049;
assign slice_143 = mul_134[17:0];
assign addW_4806 = slice_4801 + slice_4797;
assign mul_899 = slice_897 * slice_898;
assign mul_5562 = slice_5559 * slice_5561;
assign concat_1655 = {addW_1653,slice_1654};
assign lsl_6318 = mulnw_6317 << 16;
assign addW_2411 = slice_2406 + slice_2403;
assign slice_7074 = mul_7065[17:0];
assign slice_3167 = concat_3143[31:0];
assign slice_3923 = slice_3908[7:0];
assign slice_16 = slice_13[255:128];
assign mulnw_4679 = slice_4672 * slice_4678;
assign mul_772 = slice_766 * slice_768;
assign mul_5435 = slice_5431 * slice_5434;
assign slice_1528 = addW_1527[32:16];
assign mul_6191 = slice_6188 * slice_6190;
assign slice_2284 = slice_2258[7:0];
assign slice_6947 = slice_6946[32:16];
assign slice_3040 = mul_3039[35:18];
assign mulnw_3796 = slice_3789 * slice_3795;
assign slice_4552 = slice_4531[16:8];
assign mul_645 = slice_643 * slice_644;
assign addW_5308 = add_5294 + add_5307;
assign slice_1401 = addW_1400[128:64];
assign addW_6064 = add_6050 + add_6063;
assign addW_2157 = slice_2070 + slice_1984;
assign slice_6820 = slice_6819[31:18];
assign slice_2913 = mul_2912[35:18];
assign addW_7576 = concat_7570 + subW_7575;
assign slice_3669 = mul_3668[35:18];
assign concat_4425 = {mul_4420,slice_4424};
assign addW_518 = add_504 + add_517;
assign slice_5181 = concat_5180[63:32];
assign lsl_1274 = mulnw_1273 << 16;
assign subW_5937 = subW_5936 - mul_5930;
assign slice_2030 = addW_2025[15:0];
assign mul_6693 = slice_6690 * slice_6692;
assign slice_2786 = concat_2785[63:32];
assign concat_7449 = {addW_7447,slice_7448};
assign subW_3542 = concat_3541 - concat_3481;
assign concat_4298 = {mul_4293,slice_4297};
assign slice_391 = concat_345[31:0];
assign slice_5054 = slice_5053[256:128];
assign concat_1147 = {mul_1142,slice_1146};
assign lsl_5810 = mulnw_5809 << 16;
assign mulnw_1903 = slice_1896 * slice_1902;
assign slice_6566 = mul_6565[31:16];
assign slice_2659 = slice_2639[31:0];
assign mulnw_7322 = slice_7321 * slice_7318;
assign slice_3415 = concat_3414[63:32];
assign slice_4171 = mul_4170[35:18];
assign slice_264 = mul_263[35:18];
assign slice_4927 = addW_4926[65:33];
assign slice_1020 = slice_1002[15:8];
assign addW_5683 = slice_5678 + slice_5675;
assign addW_1776 = concat_1770 + subW_1775;
assign mul_6439 = slice_6434 * slice_6438;
assign concat_2532 = {addW_2530,slice_2531};
assign slice_7195 = slice_7189[15:0];
assign mulnw_3288 = slice_3281 * slice_3287;
assign mulnw_4044 = slice_4042 * slice_4043;
assign addW_137 = slice_132 + slice_127;
assign mul_4800 = slice_4797 * slice_4799;
assign slice_893 = slice_892[31:18];
assign slice_5556 = mul_5525[15:0];
assign mul_1649 = slice_1643 * slice_1645;
assign mul_6312 = slice_6306 * slice_6308;
assign slice_2405 = addW_2400[17:0];
assign addW_7068 = slice_7063 + slice_7059;
assign addW_3161 = concat_3155 + subW_3160;
assign slice_3917 = mul_3916[31:16];
assign slice_10 = IN1[1023:512];
assign slice_4673 = slice_4668[15:8];
assign slice_766 = slice_752[7:0];
assign slice_5429 = slice_5342[63:0];
assign addW_1522 = concat_1516 + subW_1521;
assign slice_6185 = mul_6176[17:0];
assign slice_2278 = slice_2260[15:8];
assign addW_6941 = concat_6913 + addW_6940;
assign slice_3034 = addW_2993[31:0];
assign slice_3790 = slice_3769[16:8];
assign add_4546 = mulnw_4543 + mulnw_4545;
assign slice_639 = addW_638[33:18];
assign mulnw_5302 = slice_5295 * slice_5301;
assign addW_1395 = concat_1307 + subW_1394;
assign mulnw_6058 = slice_6051 * slice_6057;
assign subW_2151 = subW_2150 - concat_2107;
assign concat_6814 = {addW_6812,slice_6813};
assign slice_2907 = slice_2906[63:32];
assign concat_7570 = {mul_7565,slice_7569};
assign slice_3663 = slice_3644[31:0];
assign slice_4419 = slice_4418[32:16];
assign mulnw_512 = slice_505 * slice_511;
assign mul_5175 = addW_5173 * addW_5174;
assign mul_1268 = slice_1266 * slice_1267;
assign slice_5931 = mul_5930[35:18];
assign concat_2024 = {concat_2004,slice_2023};
assign slice_6687 = concat_6686[65:33];
assign mul_2780 = addW_2778 * addW_2779;
assign addW_7443 = slice_7438 + slice_7435;
assign add_3536 = lsl_3534 + mul_3535;
assign slice_4292 = slice_4291[31:18];
assign addW_385 = concat_357 + addW_384;
assign slice_5048 = concat_5047[1023:512];
assign slice_1141 = slice_1140[31:18];
assign mul_5804 = slice_5798 * slice_5800;
assign slice_1897 = slice_1876[16:8];
assign addW_6560 = slice_6540 + slice_6522;
assign mul_2653 = addW_2651 * addW_2652;
assign concat_7316 = {mul_7311,slice_7315};
assign mul_3409 = addW_3407 * addW_3408;
assign addW_4165 = slice_4123 + slice_4083;
assign slice_258 = addW_217[31:0];
assign addW_4921 = concat_4900 + subW_4920;
assign mulnw_1014 = slice_1007 * slice_1013;
assign slice_5677 = addW_5672[17:0];
assign concat_1770 = {mul_1765,slice_1769};
assign slice_6433 = slice_6432[64:32];
assign slice_2526 = mul_2517[17:0];
assign slice_7189 = addW_7188[65:33];
assign slice_3282 = slice_3261[16:8];
assign slice_4038 = addW_4034[15:0];
assign mul_131 = slice_127 * slice_130;
assign slice_4794 = mul_4763[15:0];
assign subW_887 = mul_886 - mul_878;
assign lsl_5550 = add_5549 << 8;
assign slice_1643 = slice_1621[7:0];
assign slice_6306 = slice_6293[7:0];
assign concat_2399 = {concat_2379,slice_2398};
assign mul_7062 = slice_7059 * slice_7061;
assign concat_3155 = {mul_3150,slice_3154};
assign slice_3911 = slice_3910[64:32];
assign slice_4667 = slice_4661[15:0];
assign slice_760 = mul_759[31:16];
assign concat_5423 = {addW_5421,slice_5422};
assign concat_1516 = {mul_1511,slice_1515};
assign addW_6179 = slice_6174 + slice_6168;
assign mulnw_2272 = slice_2265 * slice_2271;
assign add_6935 = mulnw_6932 + mulnw_6934;
assign addW_3028 = add_3014 + add_3027;
assign add_3784 = mulnw_3781 + mulnw_3783;
assign mulnw_4540 = slice_4538 * slice_4539;
assign addW_633 = concat_627 + subW_632;
assign slice_5296 = slice_5275[16:8];
assign subW_1389 = subW_1388 - concat_1367;
assign slice_6052 = slice_6031[16:8];
assign add_2145 = lsl_2136 + add_2144;
assign slice_6808 = mul_6799[17:0];
assign slice_2901 = concat_2855[31:0];
assign slice_7564 = addW_7563[33:18];
assign subW_3657 = subW_3656 - mul_3650;
assign addW_4413 = concat_4385 + addW_4412;
assign slice_506 = slice_485[16:8];
assign slice_5169 = slice_5165[17:0];
assign slice_1262 = addW_1261[32:16];
assign slice_5925 = slice_5906[31:0];
assign subW_2018 = mul_2017 - mul_2009;
assign add_6681 = lsl_6679 + mul_6680;
assign slice_2774 = slice_2770[17:0];
assign slice_7437 = slice_7432[17:0];
assign mulnw_3530 = slice_3529 * slice_3526;
assign concat_4286 = {addW_4284,slice_4285};
assign add_379 = mulnw_376 + mulnw_378;
assign concat_5042 = {addW_5040,slice_5041};
assign slice_1135 = slice_1134[127:64];
assign slice_5798 = slice_5784[7:0];
assign add_1891 = mulnw_1888 + mulnw_1890;
assign slice_6554 = mul_6545[17:0];
assign slice_2647 = slice_2643[17:0];
assign slice_7310 = slice_7309[32:16];
assign slice_3403 = slice_3399[17:0];
assign slice_4159 = mul_4128[15:0];
assign addW_252 = add_238 + add_251;
assign subW_4915 = subW_4914 - mul_4908;
assign slice_1008 = slice_1003[15:8];
assign concat_5671 = {concat_5651,slice_5670};
assign slice_1764 = addW_1763[33:18];
assign slice_6427 = concat_6336[63:0];
assign addW_2520 = slice_2515 + slice_2511;
assign addW_7183 = concat_7140 + subW_7182;
assign add_3276 = mulnw_3273 + mulnw_3275;
assign addW_4032 = slice_4012 + slice_3993;
assign slice_125 = slice_16[63:0];
assign lsl_4788 = add_4787 << 8;
assign mul_881 = slice_879 * slice_880;
assign lsl_5544 = mulnw_5543 << 16;
assign add_1637 = lsl_1635 + mul_1636;
assign slice_6300 = mul_6299[31:16];
assign subW_2393 = mul_2392 - mul_2384;
assign slice_7056 = mul_7025[15:0];
assign slice_3149 = addW_3148[33:18];
assign addW_3905 = slice_3639 + slice_3374;
assign slice_4661 = addW_4660[64:32];
assign slice_754 = addW_753[65:33];
assign mul_5417 = slice_5411 * slice_5413;
assign slice_1510 = slice_1509[31:18];
assign mul_6173 = slice_6168 * slice_6172;
assign slice_2266 = slice_2261[15:8];
assign mulnw_6929 = slice_6927 * slice_6928;
assign mulnw_3022 = slice_3015 * slice_3021;
assign mulnw_3778 = slice_3776 * slice_3777;
assign slice_4534 = addW_4530[15:0];
assign concat_627 = {mul_622,slice_626};
assign add_5290 = mulnw_5287 + mulnw_5289;
assign subW_1383 = mul_1382 - mul_1374;
assign add_6046 = mulnw_6043 + mulnw_6045;
assign slice_2139 = slice_2113[7:0];
assign addW_6802 = slice_6797 + slice_6793;
assign addW_2895 = concat_2867 + addW_2894;
assign concat_7558 = {addW_7556,slice_7557};
assign slice_3651 = mul_3650[35:18];
assign add_4407 = mulnw_4404 + mulnw_4406;
assign add_500 = mulnw_497 + mulnw_499;
assign slice_5163 = slice_5143[31:0];
assign addW_1256 = concat_1250 + subW_1255;
assign subW_5919 = subW_5918 - mul_5912;
assign mul_2012 = slice_2010 * slice_2011;
assign mulnw_6675 = slice_6674 * slice_6671;
assign slice_2768 = addW_2726[31:0];
assign concat_7431 = {addW_7429,slice_7430};
assign add_3524 = lsl_3515 + add_3523;
assign slice_4280 = mul_4271[17:0];
assign mulnw_373 = slice_371 * slice_372;
assign slice_5036 = concat_4923[64:0];
assign subW_1129 = concat_1128 - concat_956;
assign slice_5792 = mul_5791[31:16];
assign mulnw_1885 = slice_1883 * slice_1884;
assign addW_6548 = slice_6543 + slice_6539;
assign slice_2641 = slice_2640[31:18];
assign slice_7304 = addW_7303[129:65];
assign slice_3397 = slice_3375[31:0];
assign lsl_4153 = add_4152 << 8;
assign mulnw_246 = slice_239 * slice_245;
assign slice_4909 = mul_4908[35:18];
assign slice_1002 = addW_997[15:0];
assign subW_5665 = mul_5664 - mul_5656;
assign concat_1758 = {addW_1756,slice_1757};
assign addW_6421 = concat_6400 + subW_6420;
assign mul_2514 = slice_2511 * slice_2513;
assign addW_7177 = add_7163 + add_7176;
assign mulnw_3270 = slice_3268 * slice_3269;
assign subW_4026 = subW_4025 - mul_4019;
assign concat_119 = {addW_117,slice_118};
assign lsl_4782 = mulnw_4781 << 16;
assign slice_875 = slice_874[127:64];
assign mul_5538 = slice_5532 * slice_5534;
assign mulnw_1631 = slice_1630 * slice_1627;
assign addW_6294 = slice_6274 + slice_6256;
assign mul_2387 = slice_2385 * slice_2386;
assign lsl_7050 = add_7049 << 8;
assign concat_3143 = {addW_3141,slice_3142};
assign subW_3899 = subW_3898 - concat_3810;
assign addW_4655 = concat_4612 + subW_4654;
assign slice_5411 = slice_5389[7:0];
assign addW_1504 = concat_1498 + subW_1503;
assign slice_6167 = slice_6166[63:32];
assign slice_2260 = slice_2253[15:0];
assign lsl_6923 = add_6922 << 8;
assign slice_3016 = slice_2995[16:8];
assign slice_3772 = addW_3768[15:0];
assign addW_4528 = slice_4508 + slice_4488;
assign slice_621 = slice_620[31:18];
assign mulnw_5284 = slice_5282 * slice_5283;
assign mul_1377 = slice_1375 * slice_1376;
assign mulnw_6040 = slice_6038 * slice_6039;
assign slice_2133 = slice_2115[15:8];
assign mul_6796 = slice_6793 * slice_6795;
assign add_2889 = mulnw_2886 + mulnw_2888;
assign mul_7552 = slice_7546 * slice_7548;
assign slice_3645 = slice_3644[63:32];
assign mulnw_4401 = slice_4399 * slice_4400;
assign mulnw_494 = slice_492 * slice_493;
assign mul_5157 = addW_5155 * addW_5156;
assign concat_1250 = {mul_1245,slice_1249};
assign slice_5913 = mul_5912[35:18];
assign slice_2006 = slice_2005[31:18];
assign add_6669 = lsl_6660 + add_6668;
assign add_2762 = lsl_2760 + mul_2761;
assign mul_7425 = slice_7419 * slice_7421;
assign slice_3518 = slice_3508[7:0];
assign addW_4274 = slice_4269 + slice_4265;
assign lsl_367 = add_366 << 8;
assign addW_5030 = concat_5009 + subW_5029;
assign concat_1123 = {addW_1121,slice_1122};
assign slice_5786 = addW_5785[65:33];
assign slice_1879 = slice_1875[15:0];
assign mul_6542 = slice_6539 * slice_6541;
assign subW_2635 = subW_2634 - concat_2591;
assign slice_7298 = concat_7185[63:0];
assign mul_3391 = addW_3389 * addW_3390;
assign lsl_4147 = mulnw_4146 << 16;
assign slice_240 = slice_219[16:8];
assign addW_4903 = slice_4883 + slice_4843;
assign concat_996 = {concat_976,slice_995};
assign mul_5659 = slice_5657 * slice_5658;
assign addW_1752 = slice_1747 + slice_1744;
assign subW_6415 = subW_6414 - mul_6408;
assign slice_2508 = concat_2507[65:33];
assign mulnw_7171 = slice_7164 * slice_7170;
assign slice_3264 = slice_3260[15:0];
assign slice_4020 = mul_4019[35:18];
assign mul_113 = slice_107 * slice_109;
assign mul_4776 = slice_4770 * slice_4772;
assign slice_869 = slice_868[255:128];
assign slice_5532 = slice_5518[7:0];
assign concat_1625 = {mul_1620,slice_1624};
assign slice_6288 = mul_6279[17:0];
assign slice_2381 = slice_2380[31:18];
assign lsl_7044 = mulnw_7043 << 16;
assign addW_3137 = slice_3132 + slice_3129;
assign subW_3893 = concat_3892 - concat_3854;
assign addW_4649 = add_4635 + add_4648;
assign subW_742 = subW_741 - concat_698;
assign add_5405 = lsl_5403 + mul_5404;
assign concat_1498 = {mul_1493,slice_1497};
assign subW_6161 = subW_6160 - concat_6072;
assign slice_2254 = slice_2253[32:16];
assign lsl_6917 = mulnw_6916 << 16;
assign add_3010 = mulnw_3007 + mulnw_3009;
assign addW_3766 = slice_3746 + slice_3727;
assign subW_4522 = subW_4521 - mul_4515;
assign addW_615 = concat_587 + addW_614;
assign slice_5278 = slice_5274[15:0];
assign slice_1371 = addW_1370[33:18];
assign slice_6034 = addW_6030[15:0];
assign mulnw_2127 = slice_2120 * slice_2126;
assign slice_6790 = concat_6789[63:32];
assign mulnw_2883 = slice_2881 * slice_2882;
assign slice_7546 = slice_7524[7:0];
assign slice_3639 = slice_3373[127:0];
assign lsl_4395 = add_4394 << 8;
assign slice_488 = slice_484[15:0];
assign slice_5151 = slice_5147[17:0];
assign slice_1244 = slice_1243[31:18];
assign slice_5907 = slice_5906[63:32];
assign subW_2000 = mul_1999 - mul_1991;
assign slice_6663 = slice_6653[7:0];
assign mulnw_2756 = slice_2755 * slice_2752;
assign slice_7419 = slice_7397[7:0];
assign slice_3512 = slice_3503[16:8];
assign mul_4268 = slice_4265 * slice_4267;
assign lsl_361 = mulnw_360 << 16;
assign subW_5024 = subW_5023 - mul_5017;
assign addW_1117 = slice_1112 + slice_1109;
assign slice_5780 = concat_5779[129:65];
assign slice_1873 = slice_1872[32:16];
assign slice_6536 = mul_6527[17:0];
assign add_2629 = lsl_2620 + add_2628;
assign addW_7292 = concat_7271 + subW_7291;
assign slice_3385 = slice_3381[17:0];
assign mul_4141 = slice_4135 * slice_4137;
assign add_234 = mulnw_231 + mulnw_233;
assign slice_4897 = mul_4888[17:0];
assign subW_990 = mul_989 - mul_981;
assign slice_5653 = slice_5652[31:18];
assign slice_1746 = slice_1741[17:0];
assign slice_6409 = mul_6408[35:18];
assign add_2502 = lsl_2500 + mul_2501;
assign slice_7165 = slice_7144[16:8];
assign slice_3258 = slice_3257[32:16];
assign slice_4014 = slice_3995[31:0];
assign slice_107 = slice_82[7:0];
assign slice_4770 = slice_4755[7:0];
assign subW_863 = concat_862 - concat_305;
assign slice_5526 = mul_5525[31:16];
assign slice_1619 = slice_1618[32:16];
assign addW_6282 = slice_6277 + slice_6273;
assign add_2375 = lsl_2366 + add_2374;
assign mul_7038 = slice_7032 * slice_7034;
assign slice_3131 = slice_3126[17:0];
assign mul_3887 = addW_3885 * addW_3886;
assign mulnw_4643 = slice_4636 * slice_4642;
assign add_736 = lsl_727 + add_735;
assign mulnw_5399 = slice_5398 * slice_5395;
assign slice_1492 = slice_1491[31:18];
assign subW_6155 = concat_6154 - concat_6116;
assign concat_2248 = {concat_1982,slice_2247};
assign mul_6911 = slice_6909 * slice_6910;
assign mulnw_3004 = slice_3002 * slice_3003;
assign subW_3760 = subW_3759 - mul_3753;
assign slice_4516 = mul_4515[35:18];
assign add_609 = mulnw_606 + mulnw_608;
assign slice_5272 = addW_5230[32:0];
assign addW_1365 = concat_1359 + subW_1364;
assign addW_6028 = slice_6008 + slice_5989;
assign slice_2121 = slice_2116[15:8];
assign mul_6784 = addW_6782 * addW_6783;
assign lsl_2877 = add_2876 << 8;
assign add_7540 = lsl_7538 + mul_7539;
assign concat_3633 = {addW_3631,slice_3632};
assign lsl_4389 = mulnw_4388 << 16;
assign slice_482 = slice_481[32:16];
assign slice_5145 = slice_5144[31:18];
assign addW_1238 = concat_1232 + subW_1237;
assign slice_5901 = slice_5900[127:64];
assign mul_1994 = slice_1992 * slice_1993;
assign slice_6657 = slice_6648[16:8];
assign add_2750 = lsl_2741 + add_2749;
assign add_7413 = lsl_7411 + mul_7412;
assign mul_3506 = slice_3503 * slice_3505;
assign slice_4262 = concat_4261[63:32];
assign mul_355 = slice_353 * slice_354;
assign slice_5018 = mul_5017[35:18];
assign slice_1111 = addW_1106[17:0];
assign concat_5774 = {addW_5772,slice_5773};
assign slice_1867 = concat_1821[31:0];
assign addW_6530 = slice_6525 + slice_6520;
assign slice_2623 = slice_2597[7:0];
assign subW_7286 = subW_7285 - mul_7279;
assign slice_3379 = slice_3378[255:128];
assign slice_4135 = slice_4122[7:0];
assign mulnw_228 = slice_226 * slice_227;
assign addW_4891 = slice_4886 + slice_4882;
assign mul_984 = slice_982 * slice_983;
assign add_5647 = lsl_5638 + add_5646;
assign concat_1740 = {addW_1738,slice_1739};
assign addW_6403 = slice_6383 + slice_6343;
assign mulnw_2496 = slice_2495 * slice_2492;
assign add_7159 = mulnw_7156 + mulnw_7158;
assign slice_3252 = concat_3206[31:0];
assign subW_4008 = subW_4007 - mul_4001;
assign add_101 = lsl_99 + mul_100;
assign slice_4764 = mul_4763[31:16];
assign concat_857 = {addW_855,slice_856};
assign slice_5520 = addW_5519[64:32];
assign addW_1613 = concat_1585 + addW_1612;
assign mul_6276 = slice_6273 * slice_6275;
assign slice_2369 = slice_2343[7:0];
assign slice_7032 = slice_7017[7:0];
assign concat_3125 = {addW_3123,slice_3124};
assign slice_3881 = addW_3877[17:0];
assign slice_4637 = slice_4616[16:8];
assign slice_730 = slice_704[7:0];
assign concat_5393 = {mul_5388,slice_5392};
assign concat_1486 = {addW_1484,slice_1485};
assign mul_6149 = addW_6147 * addW_6148;
assign subW_2242 = concat_2241 - concat_2069;
assign addW_6905 = slice_6818 + slice_6733;
assign slice_2998 = slice_2994[15:0];
assign slice_3754 = mul_3753[35:18];
assign slice_4510 = slice_4491[31:0];
assign mulnw_603 = slice_601 * slice_602;
assign add_5266 = lsl_5264 + mul_5265;
assign concat_1359 = {mul_1354,slice_1358};
assign subW_6022 = subW_6021 - mul_6015;
assign slice_2115 = addW_2110[15:0];
assign slice_6778 = slice_6774[17:0];
assign lsl_2871 = mulnw_2870 << 16;
assign mulnw_7534 = slice_7533 * slice_7530;
assign slice_3627 = mul_3618[17:0];
assign mul_4383 = slice_4381 * slice_4382;
assign slice_476 = concat_430[31:0];
assign subW_5139 = subW_5138 - concat_5117;
assign concat_1232 = {mul_1227,slice_1231};
assign subW_5895 = subW_5894 - concat_5605;
assign slice_1988 = slice_1987[127:64];
assign mul_6651 = slice_6648 * slice_6650;
assign slice_2744 = slice_2734[7:0];
assign mulnw_7407 = slice_7406 * slice_7403;
assign slice_3500 = concat_3499[63:32];
assign mul_4256 = addW_4254 * addW_4255;
assign slice_349 = addW_348[32:16];
assign addW_5012 = slice_4970 + slice_4930;
assign concat_1105 = {concat_1085,slice_1104};
assign addW_5768 = slice_5763 + slice_5760;
assign addW_1861 = concat_1833 + addW_1860;
assign mul_6524 = slice_6520 * slice_6523;
assign slice_2617 = slice_2599[15:8];
assign slice_7280 = mul_7279[35:18];
assign slice_3373 = slice_2548[255:0];
assign slice_4129 = mul_4128[31:16];
assign slice_222 = slice_218[15:0];
assign mul_4885 = slice_4882 * slice_4884;
assign slice_978 = slice_977[31:18];
assign slice_5641 = slice_5615[7:0];
assign mul_1734 = slice_1728 * slice_1730;
assign slice_6397 = mul_6388[17:0];
assign add_2490 = lsl_2481 + add_2489;
assign mulnw_7153 = slice_7151 * slice_7152;
assign addW_3246 = concat_3218 + addW_3245;
assign slice_4002 = mul_4001[35:18];
assign mulnw_95 = slice_94 * slice_90;
assign slice_4758 = slice_4757[64:32];
assign slice_851 = mul_842[17:0];
assign slice_5514 = concat_5513[127:64];
assign add_1607 = mulnw_1604 + mulnw_1606;
assign slice_6270 = mul_6261[17:0];
assign slice_2363 = slice_2345[15:8];
assign slice_7026 = mul_7025[31:16];
assign mul_3119 = slice_3113 * slice_3115;
assign addW_3875 = slice_3855 + slice_3814;
assign add_4631 = mulnw_4628 + mulnw_4630;
assign slice_724 = slice_706[15:8];
assign slice_5387 = addW_5386[32:16];
assign slice_1480 = mul_1471[17:0];
assign slice_6143 = addW_6139[17:0];
assign concat_2236 = {addW_2234,slice_2235};
assign concat_6899 = {addW_6897,slice_6898};
assign slice_2992 = slice_2991[32:16];
assign slice_3748 = slice_3729[31:0];
assign subW_4504 = subW_4503 - mul_4497;
assign lsl_597 = add_596 << 8;
assign mulnw_5260 = slice_5259 * slice_5256;
assign slice_1353 = slice_1352[31:18];
assign slice_6016 = mul_6015[35:18];
assign concat_2109 = {concat_2089,slice_2108};
assign slice_6772 = slice_6728[31:0];
assign mul_2865 = slice_2863 * slice_2864;
assign concat_7528 = {mul_7523,slice_7527};
assign addW_3621 = slice_3616 + slice_3612;
assign addW_4377 = slice_4290 + slice_4205;
assign addW_470 = concat_442 + addW_469;
assign subW_5133 = mul_5132 - mul_5124;
assign slice_1226 = slice_1225[31:18];
assign subW_5889 = concat_5888 - concat_5694;
assign concat_1982 = {addW_1980,slice_1981};
assign slice_6645 = mul_6614[15:0];
assign slice_2738 = slice_2728[16:8];
assign concat_7401 = {mul_7396,slice_7400};
assign mul_3494 = addW_3492 * addW_3493;
assign slice_4250 = slice_4246[17:0];
assign addW_343 = concat_337 + subW_342;
assign slice_5006 = mul_4975[15:0];
assign subW_1099 = mul_1098 - mul_1090;
assign slice_5762 = addW_5757[17:0];
assign add_1855 = mulnw_1852 + mulnw_1854;
assign slice_6518 = addW_6431[63:0];
assign mulnw_2611 = slice_2604 * slice_2610;
assign addW_7274 = slice_7232 + slice_7192;
assign concat_3367 = {addW_3365,slice_3366};
assign slice_4123 = addW_4082[32:0];
assign slice_216 = slice_215[32:16];
assign slice_4879 = mul_4848[15:0];
assign subW_972 = mul_971 - mul_963;
assign slice_5635 = slice_5617[15:8];
assign slice_1728 = slice_1706[7:0];
assign addW_6391 = slice_6386 + slice_6382;
assign slice_2484 = slice_2474[7:0];
assign slice_7147 = addW_7143[15:0];
assign add_3240 = mulnw_3237 + mulnw_3239;
assign slice_3996 = slice_3995[63:32];
assign slice_89 = slice_77[16:8];
assign addW_4752 = slice_4486 + slice_4199;
assign addW_845 = slice_840 + slice_836;
assign concat_5508 = {addW_5506,slice_5507};
assign mulnw_1601 = slice_1599 * slice_1600;
assign addW_6264 = slice_6259 + slice_6254;
assign mulnw_2357 = slice_2350 * slice_2356;
assign slice_7020 = slice_7019[64:32];
assign slice_3113 = slice_3091[7:0];
assign subW_3869 = subW_3868 - mul_3862;
assign mulnw_4625 = slice_4623 * slice_4624;
assign mulnw_718 = slice_711 * slice_717;
assign concat_5381 = {addW_5379,slice_5380};
assign addW_1474 = slice_1469 + slice_1465;
assign addW_6137 = slice_6117 + slice_6076;
assign addW_2230 = slice_2225 + slice_2222;
assign slice_6893 = mul_6862[15:0];
assign slice_2986 = concat_2940[31:0];
assign subW_3742 = subW_3741 - mul_3735;
assign slice_4498 = mul_4497[35:18];
assign lsl_591 = mulnw_590 << 16;
assign add_5254 = lsl_5245 + add_5253;
assign addW_1347 = concat_1319 + addW_1346;
assign slice_6010 = slice_5991[31:0];
assign subW_2103 = mul_2102 - mul_2094;
assign add_6766 = lsl_6764 + mul_6765;
assign slice_2859 = addW_2858[32:16];
assign slice_7522 = slice_7521[32:16];
assign mul_3615 = slice_3612 * slice_3614;
assign concat_4371 = {addW_4369,slice_4370};
assign add_464 = mulnw_461 + mulnw_463;
assign mul_5127 = slice_5125 * slice_5126;
assign concat_1220 = {addW_1218,slice_1219};
assign concat_5883 = {addW_5881,slice_5882};
assign slice_1976 = concat_1952[32:0];
assign lsl_6639 = add_6638 << 8;
assign mul_2732 = slice_2728 * slice_2731;
assign slice_7395 = slice_7394[32:16];
assign slice_3488 = slice_3484[17:0];
assign slice_4244 = slice_4200[31:0];
assign concat_337 = {mul_332,slice_336};
assign lsl_5000 = add_4999 << 8;
assign mul_1093 = slice_1091 * slice_1092;
assign concat_5756 = {concat_5736,slice_5755};
assign mulnw_1849 = slice_1847 * slice_1848;
assign concat_6512 = {addW_6510,slice_6511};
assign slice_2605 = slice_2600[15:8];
assign slice_7268 = mul_7237[15:0];
assign slice_3361 = concat_3337[32:0];
assign addW_4117 = add_4103 + add_4116;
assign slice_210 = concat_209[127:64];
assign lsl_4873 = add_4872 << 8;
assign mul_966 = slice_964 * slice_965;
assign mulnw_5629 = slice_5622 * slice_5628;
assign add_1722 = lsl_1720 + mul_1721;
assign mul_6385 = slice_6382 * slice_6384;
assign slice_2478 = slice_2469[16:8];
assign addW_7141 = slice_7121 + slice_7102;
assign mulnw_3234 = slice_3232 * slice_3233;
assign slice_3990 = concat_3966[31:0];
assign slice_83 = addW_78[15:0];
assign subW_4746 = subW_4745 - concat_4657;
assign mul_839 = slice_836 * slice_838;
assign mul_5502 = slice_5496 * slice_5498;
assign lsl_1595 = add_1594 << 8;
assign mul_6258 = slice_6254 * slice_6257;
assign slice_2351 = slice_2346[15:8];
assign slice_7014 = addW_6726[128:0];
assign add_3107 = lsl_3105 + mul_3106;
assign slice_3863 = mul_3862[35:18];
assign slice_4619 = addW_4615[15:0];
assign slice_712 = slice_707[15:8];
assign addW_5375 = slice_5370 + slice_5367;
assign mul_1468 = slice_1465 * slice_1467;
assign subW_6131 = subW_6130 - mul_6124;
assign slice_2224 = addW_2219[17:0];
assign lsl_6887 = add_6886 << 8;
assign addW_2980 = concat_2952 + addW_2979;
assign slice_3736 = mul_3735[35:18];
assign slice_4492 = slice_4491[63:32];
assign mul_585 = slice_583 * slice_584;
assign slice_5248 = slice_5238[7:0];
assign add_1341 = mulnw_1338 + mulnw_1340;
assign subW_6004 = subW_6003 - mul_5997;
assign mul_2097 = slice_2095 * slice_2096;
assign mulnw_6760 = slice_6759 * slice_6756;
assign addW_2853 = concat_2847 + subW_2852;
assign addW_7516 = concat_7488 + addW_7515;
assign slice_3609 = concat_3608[63:32];
assign slice_4365 = mul_4334[15:0];
assign mulnw_458 = slice_456 * slice_457;
assign slice_5121 = addW_5120[33:18];
assign slice_1214 = mul_1183[15:0];
assign addW_5877 = slice_5872 + slice_5869;
assign addW_1970 = concat_1964 + subW_1969;
assign lsl_6633 = mulnw_6632 << 16;
assign addW_2726 = slice_2639 + slice_2551;
assign concat_7389 = {addW_7387,slice_7388};
assign slice_3482 = slice_3462[31:0];
assign add_4238 = lsl_4236 + mul_4237;
assign slice_331 = slice_330[31:18];
assign lsl_4994 = mulnw_4993 << 16;
assign slice_1087 = slice_1086[31:18];
assign subW_5750 = mul_5749 - mul_5741;
assign lsl_1843 = add_1842 << 8;
assign addW_6506 = slice_6501 + slice_6498;
assign slice_2599 = addW_2594[15:0];
assign lsl_7262 = add_7261 << 8;
assign addW_3355 = concat_3349 + subW_3354;
assign mulnw_4111 = slice_4104 * slice_4110;
assign concat_204 = {addW_202,slice_203};
assign lsl_4867 = mulnw_4866 << 16;
assign slice_960 = slice_874[63:0];
assign slice_5623 = slice_5618[15:8];
assign mulnw_1716 = slice_1715 * slice_1712;
assign slice_6379 = mul_6348[15:0];
assign mul_2472 = slice_2469 * slice_2471;
assign subW_7135 = subW_7134 - mul_7128;
assign lsl_3228 = add_3227 << 8;
assign addW_3984 = concat_3978 + subW_3983;
assign slice_77 = addW_75[32:16];
assign subW_4740 = concat_4739 - concat_4701;
assign concat_833 = {concat_791,slice_832};
assign slice_5496 = slice_5474[7:0];
assign lsl_1589 = mulnw_1588 << 16;
assign slice_6252 = slice_6165[63:0];
assign slice_2345 = slice_2339[15:0];
assign concat_7008 = {addW_7006,slice_7007};
assign mulnw_3101 = slice_3100 * slice_3097;
assign slice_3857 = addW_3816[31:0];
assign addW_4613 = slice_4593 + slice_4574;
assign slice_706 = addW_701[15:0];
assign slice_5369 = slice_5364[17:0];
assign slice_1462 = concat_1461[63:32];
assign slice_6125 = mul_6124[35:18];
assign concat_2218 = {concat_2198,slice_2217};
assign lsl_6881 = mulnw_6880 << 16;
assign add_2974 = mulnw_2971 + mulnw_2973;
assign slice_3730 = slice_3729[63:32];
assign slice_4486 = addW_4198[127:0];
assign slice_579 = addW_578[128:64];
assign slice_5242 = slice_5232[16:8];
assign mulnw_1335 = slice_1333 * slice_1334;
assign slice_5998 = mul_5997[35:18];
assign slice_2091 = slice_2090[31:18];
assign add_6754 = lsl_6745 + add_6753;
assign concat_2847 = {mul_2842,slice_2846};
assign add_7510 = mulnw_7507 + mulnw_7509;
assign mul_3603 = addW_3601 * addW_3602;
assign lsl_4359 = add_4358 << 8;
assign lsl_452 = add_451 << 8;
assign addW_5115 = concat_5109 + subW_5114;
assign lsl_1208 = add_1207 << 8;
assign slice_5871 = addW_5866[17:0];
assign concat_1964 = {mul_1959,slice_1963};
assign mul_6627 = slice_6621 * slice_6623;
assign subW_2720 = subW_2719 - concat_2676;
assign slice_7383 = mul_7374[17:0];
assign mul_3476 = addW_3474 * addW_3475;
assign mulnw_4232 = slice_4231 * slice_4228;
assign addW_325 = concat_319 + subW_324;
assign mul_4988 = slice_4982 * slice_4984;
assign add_1081 = lsl_1072 + add_1080;
assign mul_5744 = slice_5742 * slice_5743;
assign lsl_1837 = mulnw_1836 << 16;
assign slice_6500 = addW_6495[17:0];
assign concat_2593 = {concat_2573,slice_2592};
assign lsl_7256 = mulnw_7255 << 16;
assign concat_3349 = {mul_3344,slice_3348};
assign slice_4105 = slice_4084[16:8];
assign mul_198 = slice_192 * slice_194;
assign mul_4861 = slice_4855 * slice_4857;
assign addW_954 = concat_911 + subW_953;
assign slice_5617 = slice_5610[15:0];
assign concat_1710 = {mul_1705,slice_1709};
assign lsl_6373 = add_6372 << 8;
assign slice_2466 = mul_2435[15:0];
assign slice_7129 = mul_7128[35:18];
assign lsl_3222 = mulnw_3221 << 16;
assign concat_3978 = {mul_3973,slice_3977};
assign concat_71 = {concat_51,slice_70};
assign mul_4734 = addW_4732 * addW_4733;
assign add_827 = lsl_818 + add_826;
assign add_5490 = lsl_5488 + mul_5489;
assign mul_1583 = slice_1581 * slice_1582;
assign concat_6246 = {addW_6244,slice_6245};
assign slice_2339 = slice_2338[64:32];
assign slice_7002 = mul_6993[17:0];
assign concat_3095 = {mul_3090,slice_3094};
assign addW_3851 = add_3837 + add_3850;
assign subW_4607 = subW_4606 - mul_4600;
assign concat_700 = {concat_680,slice_699};
assign concat_5363 = {addW_5361,slice_5362};
assign mul_1456 = addW_1454 * addW_1455;
assign slice_6119 = addW_6078[31:0];
assign subW_2212 = mul_2211 - mul_2203;
assign mul_6875 = slice_6869 * slice_6871;
assign mulnw_2968 = slice_2966 * slice_2967;
assign slice_3724 = concat_3678[31:0];
assign concat_4480 = {addW_4478,slice_4479};
assign mul_5236 = slice_5232 * slice_5235;
assign lsl_1329 = add_1328 << 8;
assign slice_5992 = slice_5991[63:32];
assign subW_2085 = mul_2084 - mul_2076;
assign slice_6748 = slice_6738[7:0];
assign slice_2841 = slice_2840[31:18];
assign mulnw_7504 = slice_7502 * slice_7503;
assign slice_3597 = slice_3593[17:0];
assign lsl_4353 = mulnw_4352 << 16;
assign lsl_446 = mulnw_445 << 16;
assign concat_5109 = {mul_5104,slice_5108};
assign lsl_1202 = mulnw_1201 << 16;
assign concat_5865 = {concat_5823,slice_5864};
assign slice_1958 = addW_1957[33:18];
assign slice_6621 = slice_6607[7:0];
assign add_2714 = lsl_2705 + add_2713;
assign addW_7377 = slice_7372 + slice_7368;
assign slice_3470 = slice_3466[17:0];
assign add_4226 = lsl_4217 + add_4225;
assign concat_319 = {mul_314,slice_318};
assign slice_4982 = slice_4969[7:0];
assign slice_1075 = slice_1049[7:0];
assign slice_5738 = slice_5737[31:18];
assign mul_1831 = slice_1829 * slice_1830;
assign concat_6494 = {concat_6474,slice_6493};
assign subW_2587 = mul_2586 - mul_2578;
assign mul_7250 = slice_7244 * slice_7246;
assign slice_3343 = addW_3342[33:18];
assign add_4099 = mulnw_4096 + mulnw_4098;
assign slice_192 = slice_170[7:0];
assign slice_4855 = slice_4841[7:0];
assign addW_948 = add_934 + add_947;
assign slice_5611 = slice_5610[32:16];
assign slice_1704 = slice_1703[32:16];
assign lsl_6367 = mulnw_6366 << 16;
assign lsl_2460 = add_2459 << 8;
assign slice_7123 = slice_7104[31:0];
assign mul_3216 = slice_3214 * slice_3215;
assign slice_3972 = addW_3971[33:18];
assign subW_65 = mul_64 - mul_56;
assign slice_4728 = addW_4724[17:0];
assign slice_821 = slice_795[7:0];
assign mulnw_5484 = slice_5483 * slice_5480;
assign addW_1577 = slice_1490 + slice_1405;
assign mul_6240 = slice_6234 * slice_6236;
assign subW_2333 = concat_2332 - concat_2294;
assign addW_6996 = slice_6991 + slice_6987;
assign slice_3089 = slice_3088[32:16];
assign mulnw_3845 = slice_3838 * slice_3844;
assign slice_4601 = mul_4600[35:18];
assign subW_694 = mul_693 - mul_685;
assign addW_5357 = slice_5352 + slice_5349;
assign slice_1450 = slice_1446[17:0];
assign addW_6113 = add_6099 + add_6112;
assign mul_2206 = slice_2204 * slice_2205;
assign slice_6869 = slice_6856[7:0];
assign lsl_2962 = add_2961 << 8;
assign addW_3718 = concat_3690 + addW_3717;
assign slice_4474 = mul_4465[17:0];
assign addW_567 = concat_479 + subW_566;
assign addW_5230 = slice_5143 + slice_5055;
assign lsl_1323 = mulnw_1322 << 16;
assign slice_5986 = concat_5940[31:0];
assign mul_2079 = slice_2077 * slice_2078;
assign slice_6742 = slice_6730[16:8];
assign addW_2835 = concat_2829 + subW_2834;
assign lsl_7498 = add_7497 << 8;
assign slice_3591 = addW_3549[31:0];
assign mul_4347 = slice_4341 * slice_4343;
assign mul_440 = slice_438 * slice_439;
assign slice_5103 = slice_5102[31:18];
assign mul_1196 = slice_1190 * slice_1192;
assign add_5859 = lsl_5850 + add_5858;
assign concat_1952 = {addW_1950,slice_1951};
assign slice_6615 = mul_6614[31:16];
assign slice_2708 = slice_2682[7:0];
assign mul_7371 = slice_7368 * slice_7370;
assign slice_3464 = slice_3463[31:18];
assign slice_4220 = slice_4210[7:0];
assign slice_313 = slice_312[31:18];
assign slice_4976 = mul_4975[31:16];
assign slice_1069 = slice_1051[15:8];
assign add_5732 = lsl_5723 + add_5731;
assign slice_1825 = addW_1824[32:16];
assign subW_6488 = mul_6487 - mul_6479;
assign mul_2581 = slice_2579 * slice_2580;
assign slice_7244 = slice_7231[7:0];
assign concat_3337 = {addW_3335,slice_3336};
assign mulnw_4093 = slice_4091 * slice_4092;
assign add_186 = lsl_184 + mul_185;
assign slice_4849 = mul_4848[31:16];
assign mulnw_942 = slice_935 * slice_941;
assign concat_5605 = {addW_5603,slice_5604};
assign slice_1698 = slice_1697[64:32];
assign mul_6361 = slice_6355 * slice_6357;
assign lsl_2454 = mulnw_2453 << 16;
assign subW_7117 = subW_7116 - mul_7110;
assign slice_3210 = addW_3209[32:16];
assign concat_3966 = {addW_3964,slice_3965};
assign mul_59 = slice_57 * slice_58;
assign addW_4722 = slice_4702 + slice_4661;
assign slice_815 = slice_797[15:8];
assign concat_5478 = {mul_5473,slice_5477};
assign concat_1571 = {addW_1569,slice_1570};
assign slice_6234 = slice_6212[7:0];
assign mul_2327 = addW_2325 * addW_2326;
assign mul_6990 = slice_6987 * slice_6989;
assign slice_3083 = addW_3082[128:64];
assign slice_3839 = slice_3818[16:8];
assign slice_4595 = slice_4576[31:0];
assign mul_688 = slice_686 * slice_687;
assign slice_5351 = slice_5344[17:0];
assign slice_1444 = slice_1401[31:0];
assign mulnw_6107 = slice_6100 * slice_6106;
assign slice_2200 = slice_2199[31:18];
assign slice_6863 = mul_6862[31:16];
assign lsl_2956 = mulnw_2955 << 16;
assign add_3712 = mulnw_3709 + mulnw_3711;
assign addW_4468 = slice_4463 + slice_4459;
assign subW_561 = subW_560 - concat_539;
assign subW_5224 = subW_5223 - concat_5180;
assign mul_1317 = slice_1315 * slice_1316;
assign addW_5980 = concat_5952 + addW_5979;
assign slice_2073 = slice_1987[63:0];
assign mul_6736 = slice_6730 * slice_6735;
assign concat_2829 = {mul_2824,slice_2828};
assign lsl_7492 = mulnw_7491 << 16;
assign add_3585 = lsl_3583 + mul_3584;
assign slice_4341 = slice_4328[7:0];
assign slice_434 = addW_433[32:16];
assign addW_5097 = concat_5069 + addW_5096;
assign slice_1190 = slice_1177[7:0];
assign slice_5853 = slice_5827[7:0];
assign mul_1946 = slice_1940 * slice_1942;
assign slice_6609 = addW_6608[65:33];
assign slice_2702 = slice_2684[15:8];
assign slice_7365 = concat_7364[63:32];
assign subW_3458 = subW_3457 - concat_3414;
assign slice_4214 = slice_4202[16:8];
assign slice_307 = slice_306[127:64];
assign slice_4970 = addW_4929[32:0];
assign mulnw_1063 = slice_1056 * slice_1062;
assign slice_5726 = slice_5700[7:0];
assign addW_1819 = concat_1813 + subW_1818;
assign mul_6482 = slice_6480 * slice_6481;
assign slice_2575 = slice_2574[31:18];
assign slice_7238 = mul_7237[31:16];
assign mul_3331 = slice_3325 * slice_3327;
assign slice_4087 = slice_4083[15:0];
assign mulnw_180 = slice_179 * slice_176;
assign slice_4843 = slice_4842[64:32];
assign slice_936 = slice_915[16:8];
assign slice_5599 = concat_5575[31:0];
assign concat_1692 = {concat_867,slice_1691};
assign slice_6355 = slice_6341[7:0];
assign mul_2448 = slice_2442 * slice_2444;
assign slice_7111 = mul_7110[35:18];
assign addW_3204 = concat_3198 + subW_3203;
assign addW_3960 = slice_3955 + slice_3952;
assign slice_53 = slice_52[31:18];
assign subW_4716 = subW_4715 - mul_4709;
assign mulnw_809 = slice_802 * slice_808;
assign slice_5472 = addW_5471[32:16];
assign slice_1565 = mul_1534[15:0];
assign add_6228 = lsl_6226 + mul_6227;
assign slice_2321 = addW_2317[17:0];
assign slice_6984 = concat_6983[65:33];
assign addW_3077 = concat_2989 + subW_3076;
assign add_3833 = mulnw_3830 + mulnw_3832;
assign subW_4589 = subW_4588 - mul_4582;
assign slice_682 = slice_681[31:18];
assign slice_5345 = slice_5344[31:18];
assign add_1438 = lsl_1436 + mul_1437;
assign slice_6101 = slice_6080[16:8];
assign add_2194 = lsl_2185 + add_2193;
assign addW_6857 = slice_6837 + slice_6819;
assign mul_2950 = slice_2948 * slice_2949;
assign mulnw_3706 = slice_3704 * slice_3705;
assign mul_4462 = slice_4459 * slice_4461;
assign subW_555 = mul_554 - mul_546;
assign add_5218 = lsl_5209 + add_5217;
assign addW_1311 = slice_1224 + slice_1139;
assign add_5974 = mulnw_5971 + mulnw_5973;
assign addW_2067 = concat_2024 + subW_2066;
assign slice_6730 = slice_6729[32:16];
assign slice_2823 = slice_2822[31:18];
assign mul_7486 = slice_7484 * slice_7485;
assign mulnw_3579 = slice_3578 * slice_3575;
assign slice_4335 = mul_4334[31:16];
assign addW_428 = concat_422 + subW_427;
assign add_5091 = mulnw_5088 + mulnw_5090;
assign slice_1184 = mul_1183[31:16];
assign slice_5847 = slice_5829[15:8];
assign slice_1940 = slice_1918[7:0];
assign slice_6603 = concat_6602[127:64];
assign mulnw_2696 = slice_2689 * slice_2695;
assign mul_7359 = addW_7357 * addW_7358;
assign add_3452 = lsl_3443 + add_3451;
assign mul_4208 = slice_4202 * slice_4207;
assign subW_301 = concat_300 - concat_124;
assign addW_4964 = add_4950 + add_4963;
assign slice_1057 = slice_1052[15:8];
assign slice_5720 = slice_5702[15:8];
assign concat_1813 = {mul_1808,slice_1812};
assign slice_6476 = slice_6475[31:18];
assign subW_2569 = mul_2568 - mul_2560;
assign slice_7232 = addW_7191[32:0];
assign slice_3325 = slice_3303[7:0];
assign slice_4081 = slice_4080[32:16];
assign concat_174 = {mul_169,slice_173};
assign slice_4837 = concat_4813[31:0];
assign add_930 = mulnw_927 + mulnw_929;
assign addW_5593 = concat_5587 + subW_5592;
assign subW_1686 = concat_1685 - concat_1133;
assign slice_6349 = mul_6348[31:16];
assign slice_2442 = slice_2428[7:0];
assign slice_7105 = slice_7104[63:32];
assign concat_3198 = {mul_3193,slice_3197};
assign slice_3954 = slice_3949[17:0];
assign subW_47 = mul_46 - mul_33;
assign slice_4710 = mul_4709[35:18];
assign slice_803 = slice_798[15:8];
assign concat_5466 = {addW_5464,slice_5465};
assign lsl_1559 = add_1558 << 8;
assign mulnw_6222 = slice_6221 * slice_6218;
assign addW_2315 = slice_2295 + slice_2253;
assign add_6978 = lsl_6976 + mul_6977;
assign subW_3071 = subW_3070 - concat_3049;
assign mulnw_3827 = slice_3825 * slice_3826;
assign slice_4583 = mul_4582[35:18];
assign subW_676 = mul_675 - mul_667;
assign addW_5339 = concat_5229 + subW_5338;
assign mulnw_1432 = slice_1431 * slice_1428;
assign add_6095 = mulnw_6092 + mulnw_6094;
assign slice_2188 = slice_2162[7:0];
assign slice_6851 = mul_6842[17:0];
assign slice_2944 = addW_2943[32:16];
assign lsl_3700 = add_3699 << 8;
assign slice_4456 = concat_4455[65:33];
assign mul_549 = slice_547 * slice_548;
assign slice_5212 = slice_5186[7:0];
assign concat_1305 = {addW_1303,slice_1304};
assign mulnw_5968 = slice_5966 * slice_5967;
assign addW_2061 = add_2047 + add_2060;
assign slice_2817 = slice_2816[127:64];
assign addW_7480 = slice_7393 + slice_7308;
assign add_3573 = lsl_3564 + add_3572;
assign addW_4329 = slice_4309 + slice_4291;
assign concat_422 = {mul_417,slice_421};
assign mulnw_5085 = slice_5083 * slice_5084;
assign addW_1178 = slice_1158 + slice_1140;
assign mulnw_5841 = slice_5834 * slice_5840;
assign add_1934 = lsl_1932 + mul_1933;
assign concat_6597 = {addW_6595,slice_6596};
assign slice_2690 = slice_2685[15:8];
assign slice_7353 = slice_7349[17:0];
assign slice_3446 = slice_3420[7:0];
assign slice_4202 = slice_4201[32:16];
assign concat_295 = {addW_293,slice_294};
assign mulnw_4958 = slice_4951 * slice_4957;
assign slice_1051 = slice_1045[15:0];
assign mulnw_5714 = slice_5707 * slice_5713;
assign slice_1807 = slice_1806[31:18];
assign add_6470 = lsl_6461 + add_6469;
assign mul_2563 = slice_2561 * slice_2562;
assign addW_7226 = add_7212 + add_7225;
assign add_3319 = lsl_3317 + mul_3318;
assign slice_4075 = concat_4029[31:0];
assign slice_168 = addW_167[32:16];
assign addW_4831 = concat_4825 + subW_4830;
assign mulnw_924 = slice_922 * slice_923;
assign concat_5587 = {mul_5582,slice_5586};
assign concat_1680 = {addW_1678,slice_1679};
assign slice_6343 = addW_6342[64:32];
assign slice_2436 = mul_2435[31:16];
assign slice_7099 = concat_7075[31:0];
assign slice_3192 = slice_3191[31:18];
assign concat_3948 = {addW_3946,slice_3947};
assign concat_41 = {mul_33,slice_40};
assign slice_4704 = addW_4663[31:0];
assign slice_797 = slice_792[15:0];
assign addW_5460 = slice_5455 + slice_5452;
assign lsl_1553 = mulnw_1552 << 16;
assign concat_6216 = {mul_6211,slice_6215};
assign subW_2309 = subW_2308 - mul_2302;
assign mulnw_6972 = slice_6971 * slice_6968;
assign subW_3065 = mul_3064 - mul_3056;
assign slice_3821 = slice_3817[15:0];
assign slice_4577 = slice_4576[63:32];
assign mul_670 = slice_668 * slice_669;
assign subW_5333 = subW_5332 - concat_5311;
assign add_1426 = lsl_1417 + add_1425;
assign mulnw_6089 = slice_6087 * slice_6088;
assign slice_2182 = slice_2164[15:8];
assign addW_6845 = slice_6840 + slice_6836;
assign addW_2938 = concat_2932 + subW_2937;
assign addW_7601 = concat_5049 + subW_7600;
assign lsl_3694 = mulnw_3693 << 16;
assign add_4450 = lsl_4448 + mul_4449;
assign slice_543 = addW_542[33:18];
assign slice_5206 = slice_5188[15:8];
assign slice_1299 = mul_1268[15:0];
assign lsl_5962 = add_5961 << 8;
assign mulnw_2055 = slice_2048 * slice_2054;
assign subW_6718 = subW_6717 - concat_6428;
assign subW_2811 = concat_2810 - concat_2638;
assign concat_7474 = {addW_7472,slice_7473};
assign slice_3567 = slice_3557[7:0];
assign slice_4323 = mul_4314[17:0];
assign slice_416 = slice_415[31:18];
assign lsl_5079 = add_5078 << 8;
assign slice_1172 = mul_1163[17:0];
assign slice_5835 = slice_5830[15:8];
assign mulnw_1928 = slice_1927 * slice_1924;
assign mul_6591 = slice_6585 * slice_6587;
assign slice_2684 = addW_2679[15:0];
assign slice_7347 = slice_7304[31:0];
assign slice_3440 = slice_3422[15:8];
assign slice_4196 = concat_4195[511:256];
assign addW_289 = slice_284 + slice_281;
assign slice_4952 = slice_4931[16:8];
assign slice_1045 = addW_1044[64:32];
assign slice_5708 = slice_5703[15:8];
assign addW_1801 = concat_1795 + subW_1800;
assign slice_6464 = slice_6438[7:0];
assign slice_2557 = slice_2556[127:64];
assign mulnw_7220 = slice_7213 * slice_7219;
assign mulnw_3313 = slice_3312 * slice_3309;
assign addW_4069 = concat_4041 + addW_4068;
assign concat_162 = {addW_160,slice_161};
assign concat_4825 = {mul_4820,slice_4824};
assign slice_918 = addW_914[15:0];
assign slice_5581 = addW_5580[33:18];
assign slice_1674 = mul_1665[17:0];
assign slice_6337 = concat_6336[127:64];
assign slice_2430 = addW_2429[65:33];
assign addW_7093 = concat_7087 + subW_7092;
assign addW_3186 = concat_3180 + subW_3185;
assign mul_3942 = slice_3936 * slice_3938;
assign addW_4698 = add_4684 + add_4697;
assign concat_791 = {addW_789,slice_790};
assign slice_5454 = slice_5449[17:0];
assign mul_1547 = slice_1541 * slice_1543;
assign slice_6210 = addW_6209[32:16];
assign slice_2303 = mul_2302[35:18];
assign add_6966 = lsl_6957 + add_6965;
assign mul_3059 = slice_3057 * slice_3058;
assign slice_3815 = slice_3814[32:16];
assign slice_4571 = concat_4525[31:0];
assign slice_664 = addW_578[63:0];
assign subW_5327 = mul_5326 - mul_5318;
assign slice_1420 = slice_1410[7:0];
assign slice_6083 = slice_6079[15:0];
assign mulnw_2176 = slice_2169 * slice_2175;
assign mul_6839 = slice_6836 * slice_6838;
assign concat_2932 = {mul_2927,slice_2931};
assign subW_7595 = subW_7594 - concat_6721;
assign mul_3688 = slice_3686 * slice_3687;
assign mulnw_4444 = slice_4443 * slice_4440;
assign addW_537 = concat_531 + subW_536;
assign mulnw_5200 = slice_5193 * slice_5199;
assign lsl_1293 = add_1292 << 8;
assign lsl_5956 = mulnw_5955 << 16;
assign slice_2049 = slice_2028[16:8];
assign subW_6712 = concat_6711 - concat_6517;
assign concat_2805 = {addW_2803,slice_2804};
assign slice_7468 = mul_7459[17:0];
assign slice_3561 = slice_3551[16:8];
assign addW_4317 = slice_4312 + slice_4308;
assign addW_410 = concat_404 + subW_409;
assign lsl_5073 = mulnw_5072 << 16;
assign addW_1166 = slice_1161 + slice_1157;
assign slice_5829 = slice_5824[15:0];
assign concat_1922 = {mul_1917,slice_1921};
assign slice_6585 = slice_6563[7:0];
assign concat_2678 = {concat_2658,slice_2677};
assign add_7341 = lsl_7339 + mul_7340;
assign mulnw_3434 = slice_3427 * slice_3433;
assign concat_4190 = {addW_4188,slice_4189};
assign slice_283 = addW_278[17:0];
assign add_4946 = mulnw_4943 + mulnw_4945;
assign addW_1039 = concat_996 + subW_1038;
assign slice_5702 = slice_5696[15:0];
assign concat_1795 = {mul_1790,slice_1794};
assign slice_6458 = slice_6440[15:8];
assign slice_2551 = slice_2550[127:64];
assign slice_7214 = slice_7193[16:8];
assign concat_3307 = {mul_3302,slice_3306};
assign add_4063 = mulnw_4060 + mulnw_4062;
assign addW_156 = slice_151 + slice_148;
assign slice_4819 = addW_4818[33:18];
assign addW_912 = slice_892 + slice_871;
assign concat_5575 = {addW_5573,slice_5574};
assign addW_1668 = slice_1663 + slice_1659;
assign concat_6331 = {addW_6329,slice_6330};
assign concat_2424 = {concat_2337,slice_2423};
assign concat_7087 = {mul_7082,slice_7086};
assign concat_3180 = {mul_3175,slice_3179};
assign slice_3936 = slice_3914[7:0];
assign slice_29 = slice_28[255:128];
assign mulnw_4692 = slice_4685 * slice_4691;
assign mul_785 = slice_779 * slice_781;
assign concat_5448 = {addW_5446,slice_5447};
assign slice_1541 = slice_1528[7:0];
assign concat_6204 = {addW_6202,slice_6203};
assign slice_2297 = slice_2256[31:0];
assign slice_6960 = slice_6950[7:0];
assign slice_3053 = addW_3052[33:18];
assign slice_3809 = concat_3763[31:0];
assign addW_4565 = concat_4537 + addW_4564;
assign addW_658 = concat_637 + subW_657;
assign mul_5321 = slice_5319 * slice_5320;
assign slice_1414 = slice_1403[16:8];
assign slice_6077 = slice_6076[32:16];
assign slice_2170 = slice_2165[15:8];
assign slice_6833 = mul_6824[17:0];
assign slice_2926 = slice_2925[31:18];
assign subW_7589 = concat_7588 - concat_7013;
assign slice_3682 = addW_3681[32:16];
assign add_4438 = lsl_4429 + add_4437;
assign concat_531 = {mul_526,slice_530};
assign slice_5194 = slice_5189[15:8];
assign lsl_1287 = mulnw_1286 << 16;
assign mul_5950 = slice_5948 * slice_5949;
assign add_2043 = mulnw_2040 + mulnw_2042;
assign concat_6706 = {addW_6704,slice_6705};
assign addW_2799 = slice_2794 + slice_2791;
assign addW_7462 = slice_7457 + slice_7453;
assign mul_3555 = slice_3551 * slice_3554;
assign mul_4311 = slice_4308 * slice_4310;
assign concat_404 = {mul_399,slice_403};
assign mul_5067 = slice_5065 * slice_5066;
assign mul_1160 = slice_1157 * slice_1159;
assign concat_5823 = {addW_5821,slice_5822};
assign slice_1916 = slice_1915[32:16];
assign add_6579 = lsl_6577 + mul_6578;
assign subW_2672 = mul_2671 - mul_2663;
assign mulnw_7335 = slice_7334 * slice_7331;
assign slice_3428 = slice_3423[15:8];
assign slice_4184 = concat_4160[32:0];
assign mulnw_4940 = slice_4938 * slice_4939;
assign addW_1033 = add_1019 + add_1032;
assign slice_5696 = slice_5695[64:32];
assign slice_1789 = slice_1788[31:18];
assign mulnw_6452 = slice_6445 * slice_6451;
assign addW_2545 = concat_1692 + subW_2544;
assign add_7208 = mulnw_7205 + mulnw_7207;
assign slice_3301 = slice_3300[32:16];
assign mulnw_4057 = slice_4055 * slice_4056;
assign slice_150 = slice_145[17:0];
assign concat_4813 = {addW_4811,slice_4812};
assign subW_906 = subW_905 - mul_899;
assign addW_5569 = slice_5564 + slice_5561;
assign mul_1662 = slice_1659 * slice_1661;
assign mul_6325 = slice_6319 * slice_6321;
assign subW_2418 = concat_2417 - concat_2379;
assign slice_7081 = addW_7080[33:18];
assign slice_3174 = slice_3173[31:18];
assign add_3930 = lsl_3928 + mul_3929;
assign slice_4686 = slice_4665[16:8];
assign slice_779 = slice_757[7:0];
assign addW_5442 = slice_5437 + slice_5434;
assign slice_1535 = mul_1534[31:16];
assign addW_6198 = slice_6193 + slice_6190;
assign addW_2291 = add_2277 + add_2290;
assign slice_6954 = slice_6945[16:8];
assign addW_3047 = concat_3041 + subW_3046;
assign addW_3803 = concat_3775 + addW_3802;
assign add_4559 = mulnw_4556 + mulnw_4558;
assign subW_652 = subW_651 - mul_645;
assign slice_5315 = addW_5314[33:18];
assign mul_1408 = slice_1403 * slice_1407;
assign slice_6071 = concat_6025[31:0];
assign slice_2164 = slice_2158[15:0];
assign addW_6827 = slice_6822 + slice_6817;
assign addW_2920 = concat_2914 + subW_2919;
assign concat_7583 = {addW_7581,slice_7582};
assign addW_3676 = concat_3670 + subW_3675;
assign slice_4432 = slice_4422[7:0];
assign slice_525 = slice_524[31:18];
assign slice_5188 = addW_5183[15:0];
assign mul_1281 = slice_1275 * slice_1277;
assign slice_5944 = addW_5943[32:16];
assign mulnw_2037 = slice_2035 * slice_2036;
assign addW_6700 = slice_6695 + slice_6692;
assign slice_2793 = addW_2788[17:0];
assign mul_7456 = slice_7453 * slice_7455;
assign addW_3549 = slice_3462 + slice_3375;
assign slice_4305 = mul_4296[17:0];
assign slice_398 = slice_397[31:18];
assign slice_5061 = slice_5060[128:64];
assign slice_1154 = mul_1145[17:0];
assign mul_5817 = slice_5811 * slice_5813;
assign addW_1910 = concat_1882 + addW_1909;
assign mulnw_6573 = slice_6572 * slice_6569;
assign mul_2666 = slice_2664 * slice_2665;
assign add_7329 = lsl_7320 + add_7328;
assign slice_3422 = addW_3417[15:0];
assign addW_4178 = concat_4172 + subW_4177;
assign addW_271 = concat_265 + subW_270;
assign slice_4934 = slice_4930[15:0];
assign mulnw_1027 = slice_1020 * slice_1026;
assign subW_5690 = concat_5689 - concat_5651;
assign concat_1783 = {addW_1781,slice_1782};
assign slice_6446 = slice_6441[15:8];
assign subW_2539 = subW_2538 - concat_2246;
assign mulnw_7202 = slice_7200 * slice_7201;
assign addW_3295 = concat_3267 + addW_3294;
assign lsl_4051 = add_4050 << 8;
assign concat_144 = {addW_142,slice_143};
assign addW_4807 = slice_4802 + slice_4799;
assign slice_900 = mul_899[35:18];
assign slice_5563 = slice_5558[17:0];
assign slice_1656 = concat_1655[65:33];
assign slice_6319 = slice_6297[7:0];
assign mul_2412 = addW_2410 * addW_2411;
assign concat_7075 = {addW_7073,slice_7074};
assign concat_3168 = {addW_3166,slice_3167};
assign mulnw_3924 = slice_3923 * slice_3920;
assign add_4680 = mulnw_4677 + mulnw_4679;
assign add_773 = lsl_771 + mul_772;
assign slice_5436 = slice_5430[17:0];
assign addW_1529 = slice_1509 + slice_1491;
assign slice_6192 = slice_6187[17:0];
assign mulnw_2285 = slice_2278 * slice_2284;
assign mul_6948 = slice_6945 * slice_6947;
assign concat_3041 = {mul_3036,slice_3040};
assign add_3797 = mulnw_3794 + mulnw_3796;
assign mulnw_4553 = slice_4551 * slice_4552;
assign slice_646 = mul_645[35:18];
assign addW_5309 = concat_5281 + addW_5308;
assign slice_1402 = slice_1401[64:32];
assign addW_6065 = concat_6037 + addW_6064;
assign slice_2158 = addW_2157[64:32];
assign mul_6821 = slice_6817 * slice_6820;
assign concat_2914 = {mul_2909,slice_2913};
assign slice_7577 = mul_7568[17:0];
assign concat_3670 = {mul_3665,slice_3669};
assign slice_4426 = slice_4417[16:8];
assign addW_519 = concat_491 + addW_518;
assign concat_5182 = {concat_5162,slice_5181};
assign slice_1275 = slice_1262[7:0];
assign addW_5938 = concat_5932 + subW_5937;
assign slice_2031 = addW_2027[15:0];
assign slice_6694 = addW_6689[17:0];
assign concat_2787 = {concat_2767,slice_2786};
assign slice_7450 = concat_7449[63:32];
assign subW_3543 = subW_3542 - concat_3499;
assign addW_4299 = slice_4294 + slice_4289;
assign concat_392 = {addW_390,slice_391};
assign slice_5055 = slice_5054[128:64];
assign addW_1148 = slice_1143 + slice_1137;
assign slice_5811 = slice_5789[7:0];
assign add_1904 = mulnw_1901 + mulnw_1903;
assign concat_6567 = {mul_6562,slice_6566};
assign slice_2660 = slice_2659[31:18];
assign slice_7323 = slice_7313[7:0];
assign concat_3416 = {concat_3396,slice_3415};
assign concat_4172 = {mul_4167,slice_4171};
assign concat_265 = {mul_260,slice_264};
assign slice_4928 = slice_4927[32:16];
assign slice_1021 = slice_1000[16:8];
assign mul_5684 = addW_5682 * addW_5683;
assign slice_1777 = mul_1768[17:0];
assign slice_6440 = slice_6433[15:0];
assign subW_2533 = concat_2532 - concat_2337;
assign slice_7196 = slice_7192[15:0];
assign add_3289 = mulnw_3286 + mulnw_3288;
assign lsl_4045 = mulnw_4044 << 16;
assign addW_138 = slice_133 + slice_130;
assign slice_4801 = slice_4796[17:0];
assign slice_894 = slice_875[31:0];
assign concat_5557 = {addW_5555,slice_5556};
assign add_1650 = lsl_1648 + mul_1649;
assign add_6313 = lsl_6311 + mul_6312;
assign slice_2406 = addW_2402[17:0];
assign addW_7069 = slice_7064 + slice_7061;
assign slice_3162 = mul_3153[17:0];
assign concat_3918 = {mul_3913,slice_3917};
assign mulnw_4674 = slice_4672 * slice_4673;
assign mulnw_767 = slice_766 * slice_763;
assign slice_5430 = slice_5429[63:32];
assign slice_1523 = mul_1514[17:0];
assign concat_6186 = {addW_6184,slice_6185};
assign slice_2279 = slice_2258[16:8];
assign slice_6942 = mul_6911[15:0];
assign slice_3035 = slice_3034[31:18];
assign mulnw_3791 = slice_3789 * slice_3790;
assign lsl_4547 = add_4546 << 8;
assign addW_640 = slice_620 + slice_580;
assign add_5303 = mulnw_5300 + mulnw_5302;
assign slice_1396 = concat_1305[63:0];
assign add_6059 = mulnw_6056 + mulnw_6058;
assign addW_2152 = concat_2109 + subW_2151;
assign slice_6815 = slice_6727[63:0];
assign slice_2908 = slice_2907[31:18];
assign addW_7571 = slice_7566 + slice_7562;
assign slice_3664 = slice_3663[31:18];
assign mul_4420 = slice_4417 * slice_4419;
assign add_513 = mulnw_510 + mulnw_512;
assign subW_5176 = mul_5175 - mul_5167;
assign slice_1269 = mul_1268[31:16];
assign concat_5932 = {mul_5927,slice_5931};
assign addW_2025 = slice_2005 + slice_1985;
assign concat_6688 = {concat_6646,slice_6687};
assign subW_2781 = mul_2780 - mul_2772;
assign mul_7444 = addW_7442 * addW_7443;
assign add_3537 = lsl_3528 + add_3536;
assign mul_4293 = slice_4289 * slice_4292;
assign slice_386 = mul_355[15:0];
assign concat_5049 = {concat_2547,slice_5048};
assign mul_1142 = slice_1137 * slice_1141;
assign add_5805 = lsl_5803 + mul_5804;
assign mulnw_1898 = slice_1896 * slice_1897;
assign slice_6561 = addW_6560[32:16];
assign subW_2654 = mul_2653 - mul_2645;
assign slice_7317 = slice_7306[16:8];
assign subW_3410 = mul_3409 - mul_3401;
assign slice_4166 = addW_4165[33:18];
assign slice_259 = slice_258[31:18];
assign slice_4922 = concat_4898[31:0];
assign add_1015 = mulnw_1012 + mulnw_1014;
assign slice_5678 = addW_5674[17:0];
assign addW_1771 = slice_1766 + slice_1762;
assign slice_6434 = slice_6433[32:16];
assign concat_2527 = {addW_2525,slice_2526};
assign slice_7190 = slice_7189[32:16];
assign mulnw_3283 = slice_3281 * slice_3282;
assign mul_4039 = slice_4037 * slice_4038;
assign slice_132 = slice_126[17:0];
assign concat_4795 = {addW_4793,slice_4794};
assign subW_888 = subW_887 - mul_881;
assign mul_5551 = slice_5545 * slice_5547;
assign mulnw_1644 = slice_1643 * slice_1640;
assign mulnw_6307 = slice_6306 * slice_6303;
assign addW_2400 = slice_2380 + slice_2339;
assign slice_7063 = slice_7058[17:0];
assign addW_3156 = slice_3151 + slice_3147;
assign slice_3912 = slice_3911[32:16];
assign slice_4668 = slice_4664[15:0];
assign concat_761 = {mul_756,slice_760};
assign subW_5424 = concat_5423 - concat_5363;
assign addW_1517 = slice_1512 + slice_1508;
assign addW_6180 = slice_6175 + slice_6172;
assign add_2273 = mulnw_2270 + mulnw_2272;
assign lsl_6936 = add_6935 << 8;
assign addW_3029 = concat_3001 + addW_3028;
assign lsl_3785 = add_3784 << 8;
assign lsl_4541 = mulnw_4540 << 16;
assign slice_634 = mul_625[17:0];
assign mulnw_5297 = slice_5295 * slice_5296;
assign addW_1390 = concat_1369 + subW_1389;
assign mulnw_6053 = slice_6051 * slice_6052;
assign addW_2146 = add_2132 + add_2145;
assign concat_6809 = {addW_6807,slice_6808};
assign concat_2902 = {addW_2900,slice_2901};
assign mul_7565 = slice_7562 * slice_7564;
assign addW_3658 = concat_3652 + subW_3657;
assign slice_4414 = mul_4383[15:0];
assign mulnw_507 = slice_505 * slice_506;
assign mul_5170 = slice_5168 * slice_5169;
assign addW_1263 = slice_1243 + slice_1225;
assign slice_5926 = slice_5925[31:18];
assign subW_2019 = subW_2018 - mul_2012;
assign add_6682 = lsl_6673 + add_6681;
assign mul_2775 = slice_2773 * slice_2774;
assign slice_7438 = slice_7434[17:0];
assign slice_3531 = slice_3505[7:0];
assign slice_4287 = slice_4199[63:0];
assign lsl_380 = add_379 << 8;
assign subW_5043 = concat_5042 - concat_3372;
assign slice_1136 = slice_1135[63:32];
assign mulnw_5799 = slice_5798 * slice_5795;
assign lsl_1892 = add_1891 << 8;
assign concat_6555 = {addW_6553,slice_6554};
assign mul_2648 = slice_2646 * slice_2647;
assign mul_7311 = slice_7306 * slice_7310;
assign mul_3404 = slice_3402 * slice_3403;
assign concat_4160 = {addW_4158,slice_4159};
assign addW_253 = concat_225 + addW_252;
assign addW_4916 = concat_4910 + subW_4915;
assign mulnw_1009 = slice_1007 * slice_1008;
assign addW_5672 = slice_5652 + slice_5610;
assign mul_1765 = slice_1762 * slice_1764;
assign concat_6428 = {addW_6426,slice_6427};
assign addW_2521 = slice_2516 + slice_2513;
assign slice_7184 = concat_7138[31:0];
assign lsl_3277 = add_3276 << 8;
assign slice_4033 = addW_4032[32:16];
assign slice_126 = slice_125[63:32];
assign mul_4789 = slice_4783 * slice_4785;
assign slice_882 = mul_881[35:18];
assign slice_5545 = slice_5523[7:0];
assign add_1638 = lsl_1629 + add_1637;
assign concat_6301 = {mul_6296,slice_6300};
assign subW_2394 = subW_2393 - mul_2387;
assign concat_7057 = {addW_7055,slice_7056};
assign mul_3150 = slice_3147 * slice_3149;
assign slice_3906 = addW_3905[128:64];
assign slice_4662 = slice_4661[32:16];
assign slice_755 = slice_754[32:16];
assign add_5418 = lsl_5416 + mul_5417;
assign mul_1511 = slice_1508 * slice_1510;
assign slice_6174 = slice_6167[17:0];
assign mulnw_2267 = slice_2265 * slice_2266;
assign lsl_6930 = mulnw_6929 << 16;
assign add_3023 = mulnw_3020 + mulnw_3022;
assign lsl_3779 = mulnw_3778 << 16;
assign mul_4535 = slice_4533 * slice_4534;
assign addW_628 = slice_623 + slice_619;
assign lsl_5291 = add_5290 << 8;
assign subW_1384 = subW_1383 - mul_1377;
assign lsl_6047 = add_6046 << 8;
assign mulnw_2140 = slice_2133 * slice_2139;
assign addW_6803 = slice_6798 + slice_6795;
assign slice_2896 = mul_2865[15:0];
assign slice_7559 = concat_7558[65:33];
assign concat_3652 = {mul_3647,slice_3651};
assign lsl_4408 = add_4407 << 8;
assign lsl_501 = add_500 << 8;
assign slice_5164 = slice_5163[31:18];
assign slice_1257 = mul_1248[17:0];
assign addW_5920 = concat_5914 + subW_5919;
assign slice_2013 = mul_2012[35:18];
assign slice_6676 = slice_6650[7:0];
assign slice_2769 = slice_2768[31:18];
assign slice_7432 = slice_7390[31:0];
assign slice_3525 = slice_3507[15:8];
assign concat_4281 = {addW_4279,slice_4280};
assign lsl_374 = mulnw_373 << 16;
assign concat_5037 = {addW_5035,slice_5036};
assign subW_1130 = subW_1129 - concat_1041;
assign concat_5793 = {mul_5788,slice_5792};
assign lsl_1886 = mulnw_1885 << 16;
assign addW_6549 = slice_6544 + slice_6541;
assign slice_2642 = slice_2556[63:0];
assign slice_7305 = slice_7304[64:32];
assign slice_3398 = slice_3397[31:18];
assign mul_4154 = slice_4148 * slice_4150;
assign add_247 = mulnw_244 + mulnw_246;
assign concat_4910 = {mul_4905,slice_4909};
assign slice_1003 = addW_999[15:0];
assign subW_5666 = subW_5665 - mul_5659;
assign slice_1759 = concat_1758[63:32];
assign slice_6422 = concat_6398[31:0];
assign slice_2515 = addW_2510[17:0];
assign addW_7178 = concat_7150 + addW_7177;
assign lsl_3271 = mulnw_3270 << 16;
assign addW_4027 = concat_4021 + subW_4026;
assign subW_120 = concat_119 - concat_51;
assign slice_4783 = slice_4761[7:0];
assign slice_876 = slice_875[63:32];
assign add_5539 = lsl_5537 + mul_5538;
assign slice_1632 = slice_1622[7:0];
assign slice_6295 = addW_6294[32:16];
assign slice_2388 = mul_2387[35:18];
assign mul_7051 = slice_7045 * slice_7047;
assign slice_3144 = concat_3143[63:32];
assign addW_3900 = concat_3812 + subW_3899;
assign slice_4656 = concat_4610[31:0];
assign mulnw_5412 = slice_5411 * slice_5408;
assign slice_1505 = mul_1496[17:0];
assign slice_6168 = slice_6167[31:18];
assign slice_2261 = slice_2257[15:0];
assign mul_6924 = slice_6918 * slice_6920;
assign mulnw_3017 = slice_3015 * slice_3016;
assign mul_3773 = slice_3771 * slice_3772;
assign slice_4529 = addW_4528[32:16];
assign mul_622 = slice_619 * slice_621;
assign lsl_5285 = mulnw_5284 << 16;
assign slice_1378 = mul_1377[35:18];
assign lsl_6041 = mulnw_6040 << 16;
assign slice_2134 = slice_2113[16:8];
assign slice_6797 = addW_6792[17:0];
assign lsl_2890 = add_2889 << 8;
assign add_7553 = lsl_7551 + mul_7552;
assign slice_3646 = slice_3645[31:18];
assign lsl_4402 = mulnw_4401 << 16;
assign lsl_495 = mulnw_494 << 16;
assign subW_5158 = mul_5157 - mul_5149;
assign addW_1251 = slice_1246 + slice_1242;
assign concat_5914 = {mul_5909,slice_5913};
assign slice_2007 = slice_1988[31:0];
assign slice_6670 = slice_6652[15:8];
assign add_2763 = lsl_2754 + add_2762;
assign add_7426 = lsl_7424 + mul_7425;
assign mulnw_3519 = slice_3512 * slice_3518;
assign addW_4275 = slice_4270 + slice_4267;
assign mul_368 = slice_362 * slice_364;
assign slice_5031 = concat_5007[32:0];
assign subW_1124 = concat_1123 - concat_1085;
assign slice_5787 = slice_5786[32:16];
assign mul_1880 = slice_1878 * slice_1879;
assign slice_6543 = slice_6538[17:0];
assign addW_2636 = concat_2593 + subW_2635;
assign concat_7299 = {addW_7297,slice_7298};
assign subW_3392 = mul_3391 - mul_3383;
assign slice_4148 = slice_4126[7:0];
assign mulnw_241 = slice_239 * slice_240;
assign slice_4904 = addW_4903[33:18];
assign addW_997 = slice_977 + slice_958;
assign slice_5660 = mul_5659[35:18];
assign mul_1753 = addW_1751 * addW_1752;
assign addW_6416 = concat_6410 + subW_6415;
assign concat_2509 = {concat_2467,slice_2508};
assign add_7172 = mulnw_7169 + mulnw_7171;
assign mul_3265 = slice_3263 * slice_3264;
assign concat_4021 = {mul_4016,slice_4020};
assign add_114 = lsl_112 + mul_113;
assign add_4777 = lsl_4775 + mul_4776;
assign slice_870 = slice_869[127:64];
assign mulnw_5533 = slice_5532 * slice_5529;
assign slice_1626 = slice_1617[16:8];
assign concat_6289 = {addW_6287,slice_6288};
assign slice_2382 = slice_2341[31:0];
assign slice_7045 = slice_7023[7:0];
assign mul_3138 = addW_3136 * addW_3137;
assign subW_3894 = subW_3893 - concat_3872;
assign addW_4650 = concat_4622 + addW_4649;
assign addW_743 = concat_700 + subW_742;
assign add_5406 = lsl_5397 + add_5405;
assign addW_1499 = slice_1494 + slice_1489;
assign addW_6162 = concat_6074 + subW_6161;
assign addW_2255 = slice_1987 + slice_1701;
assign slice_6918 = slice_6904[7:0];
assign lsl_3011 = add_3010 << 8;
assign slice_3767 = addW_3766[32:16];
assign addW_4523 = concat_4517 + subW_4522;
assign slice_616 = mul_585[15:0];
assign mul_5279 = slice_5277 * slice_5278;
assign addW_1372 = slice_1352 + slice_1312;
assign mul_6035 = slice_6033 * slice_6034;
assign add_2128 = mulnw_2125 + mulnw_2127;
assign concat_6791 = {concat_6771,slice_6790};
assign lsl_2884 = mulnw_2883 << 16;
assign mulnw_7547 = slice_7546 * slice_7543;
assign slice_3640 = slice_3639[127:64];
assign mul_4396 = slice_4390 * slice_4392;
assign mul_489 = slice_487 * slice_488;
assign mul_5152 = slice_5150 * slice_5151;
assign mul_1245 = slice_1242 * slice_1244;
assign slice_5908 = slice_5907[31:18];
assign subW_2001 = subW_2000 - mul_1994;
assign mulnw_6664 = slice_6657 * slice_6663;
assign slice_2757 = slice_2731[7:0];
assign mulnw_7420 = slice_7419 * slice_7416;
assign slice_3513 = slice_3508[15:8];
assign slice_4269 = addW_4264[17:0];
assign slice_362 = slice_349[7:0];
assign addW_5025 = concat_5019 + subW_5024;
assign mul_1118 = addW_1116 * addW_1117;
assign concat_5781 = {concat_5694,slice_5780};
assign addW_1874 = slice_1787 + slice_1702;
assign concat_6537 = {addW_6535,slice_6536};
assign addW_2630 = add_2616 + add_2629;
assign slice_7293 = concat_7269[32:0];
assign mul_3386 = slice_3384 * slice_3385;
assign add_4142 = lsl_4140 + mul_4141;
assign lsl_235 = add_234 << 8;
assign concat_4898 = {addW_4896,slice_4897};
assign subW_991 = subW_990 - mul_984;
assign slice_5654 = slice_5613[31:0];
assign slice_1747 = slice_1743[17:0];
assign concat_6410 = {mul_6405,slice_6409};
assign add_2503 = lsl_2494 + add_2502;
assign mulnw_7166 = slice_7164 * slice_7165;
assign addW_3259 = slice_3172 + slice_3087;
assign slice_4015 = slice_4014[31:18];
assign mulnw_108 = slice_107 * slice_104;
assign mulnw_4771 = slice_4770 * slice_4767;
assign subW_864 = subW_863 - concat_569;
assign concat_5527 = {mul_5522,slice_5526};
assign mul_1620 = slice_1617 * slice_1619;
assign addW_6283 = slice_6278 + slice_6275;
assign addW_2376 = add_2362 + add_2375;
assign add_7039 = lsl_7037 + mul_7038;
assign slice_3132 = slice_3128[17:0];
assign subW_3888 = mul_3887 - mul_3879;
assign add_4644 = mulnw_4641 + mulnw_4643;
assign addW_737 = add_723 + add_736;
assign slice_5400 = slice_5390[7:0];
assign mul_1493 = slice_1489 * slice_1492;
assign subW_6156 = subW_6155 - concat_6134;
assign slice_6912 = mul_6911[31:16];
assign lsl_3005 = mulnw_3004 << 16;
assign addW_3761 = concat_3755 + subW_3760;
assign concat_4517 = {mul_4512,slice_4516};
assign lsl_610 = add_609 << 8;
assign slice_5273 = slice_5272[32:16];
assign slice_1366 = mul_1357[17:0];
assign slice_6029 = addW_6028[32:16];
assign mulnw_2122 = slice_2120 * slice_2121;
assign subW_6785 = mul_6784 - mul_6776;
assign mul_2878 = slice_2872 * slice_2874;
assign add_7541 = lsl_7532 + add_7540;
assign subW_3634 = concat_3633 - concat_3461;
assign slice_4390 = slice_4376[7:0];
assign addW_483 = slice_396 + slice_311;
assign slice_5146 = slice_5060[63:0];
assign slice_1239 = mul_1230[17:0];
assign slice_5902 = slice_5901[63:32];
assign slice_1995 = mul_1994[35:18];
assign slice_6658 = slice_6653[15:8];
assign slice_2751 = slice_2733[15:8];
assign add_7414 = lsl_7405 + add_7413;
assign slice_3507 = addW_3502[15:0];
assign concat_4263 = {concat_4243,slice_4262};
assign slice_356 = mul_355[31:16];
assign concat_5019 = {mul_5014,slice_5018};
assign slice_1112 = addW_1108[17:0];
assign subW_5775 = concat_5774 - concat_5736;
assign concat_1868 = {addW_1866,slice_1867};
assign addW_6531 = slice_6526 + slice_6523;
assign mulnw_2624 = slice_2617 * slice_2623;
assign addW_7287 = concat_7281 + subW_7286;
assign slice_3380 = slice_3379[127:64];
assign mulnw_4136 = slice_4135 * slice_4132;
assign lsl_229 = mulnw_228 << 16;
assign addW_4892 = slice_4887 + slice_4884;
assign slice_985 = mul_984[35:18];
assign addW_5648 = add_5634 + add_5647;
assign slice_1741 = slice_1697[31:0];
assign slice_6404 = addW_6403[33:18];
assign slice_2497 = slice_2471[7:0];
assign lsl_7160 = add_7159 << 8;
assign concat_3253 = {addW_3251,slice_3252};
assign addW_4009 = concat_4003 + subW_4008;
assign add_102 = lsl_92 + add_101;
assign concat_4765 = {mul_4760,slice_4764};
assign subW_858 = concat_857 - concat_660;
assign slice_5521 = slice_5520[32:16];
assign slice_1614 = mul_1583[15:0];
assign slice_6277 = slice_6272[17:0];
assign mulnw_2370 = slice_2363 * slice_2369;
assign mulnw_7033 = slice_7032 * slice_7029;
assign slice_3126 = slice_3083[31:0];
assign mul_3882 = slice_3880 * slice_3881;
assign mulnw_4638 = slice_4636 * slice_4637;
assign mulnw_731 = slice_724 * slice_730;
assign slice_5394 = slice_5385[16:8];
assign slice_1487 = addW_1400[63:0];
assign subW_6150 = mul_6149 - mul_6141;
assign subW_2243 = subW_2242 - concat_2154;
assign slice_6906 = addW_6905[65:33];
assign mul_2999 = slice_2997 * slice_2998;
assign concat_3755 = {mul_3750,slice_3754};
assign slice_4511 = slice_4510[31:18];
assign lsl_604 = mulnw_603 << 16;
assign add_5267 = lsl_5258 + add_5266;
assign addW_1360 = slice_1355 + slice_1351;
assign addW_6023 = concat_6017 + subW_6022;
assign slice_2116 = addW_2112[15:0];
assign mul_6779 = slice_6777 * slice_6778;
assign slice_2872 = slice_2859[7:0];
assign slice_7535 = slice_7525[7:0];
assign concat_3628 = {addW_3626,slice_3627};
assign slice_4384 = mul_4383[31:16];
assign concat_477 = {addW_475,slice_476};
assign addW_5140 = concat_5119 + subW_5139;
assign addW_1233 = slice_1228 + slice_1223;
assign addW_5896 = concat_5607 + subW_5895;
assign slice_1989 = slice_1988[63:32];
assign slice_6652 = slice_6647[15:0];
assign mulnw_2745 = slice_2738 * slice_2744;
assign slice_7408 = slice_7398[7:0];
assign concat_3501 = {concat_3481,slice_3500};
assign subW_4257 = mul_4256 - mul_4248;
assign addW_350 = slice_330 + slice_312;
assign slice_5013 = addW_5012[33:18];
assign addW_1106 = slice_1086 + slice_1045;
assign mul_5769 = addW_5767 * addW_5768;
assign slice_1862 = mul_1831[15:0];
assign slice_6525 = slice_6519[17:0];
assign slice_2618 = slice_2597[16:8];
assign concat_7281 = {mul_7276,slice_7280};
assign slice_3374 = slice_3373[255:128];
assign concat_4130 = {mul_4125,slice_4129};
assign mul_223 = slice_221 * slice_222;
assign slice_4886 = slice_4881[17:0];
assign slice_979 = slice_960[31:0];
assign mulnw_5642 = slice_5635 * slice_5641;
assign add_1735 = lsl_1733 + mul_1734;
assign concat_6398 = {addW_6396,slice_6397};
assign slice_2491 = slice_2473[15:8];
assign lsl_7154 = mulnw_7153 << 16;
assign slice_3247 = mul_3216[15:0];
assign concat_4003 = {mul_3998,slice_4002};
assign slice_96 = slice_83[7:0];
assign slice_4759 = slice_4758[32:16];
assign concat_852 = {addW_850,slice_851};
assign concat_5515 = {concat_5428,slice_5514};
assign lsl_1608 = add_1607 << 8;
assign concat_6271 = {addW_6269,slice_6270};
assign slice_2364 = slice_2343[16:8];
assign concat_7027 = {mul_7022,slice_7026};
assign add_3120 = lsl_3118 + mul_3119;
assign slice_3876 = addW_3875[33:18];
assign lsl_4632 = add_4631 << 8;
assign slice_725 = slice_704[16:8];
assign mul_5388 = slice_5385 * slice_5387;
assign concat_1481 = {addW_1479,slice_1480};
assign mul_6144 = slice_6142 * slice_6143;
assign subW_2237 = concat_2236 - concat_2198;
assign slice_6900 = concat_6899[127:64];
assign addW_2993 = slice_2906 + slice_2821;
assign slice_3749 = slice_3748[31:18];
assign addW_4505 = concat_4499 + subW_4504;
assign mul_598 = slice_592 * slice_594;
assign slice_5261 = slice_5235[7:0];
assign mul_1354 = slice_1351 * slice_1353;
assign concat_6017 = {mul_6012,slice_6016};
assign addW_2110 = slice_2090 + slice_2071;
assign slice_6773 = slice_6772[31:18];
assign slice_2866 = mul_2865[31:16];
assign slice_7529 = slice_7520[16:8];
assign addW_3622 = slice_3617 + slice_3614;
assign slice_4378 = addW_4377[65:33];
assign slice_471 = mul_440[15:0];
assign subW_5134 = subW_5133 - mul_5127;
assign mul_1227 = slice_1223 * slice_1226;
assign subW_5890 = subW_5889 - concat_5779;
assign slice_1983 = addW_1695[127:0];
assign concat_6646 = {addW_6644,slice_6645};
assign slice_2739 = slice_2734[15:8];
assign slice_7402 = slice_7392[16:8];
assign subW_3495 = mul_3494 - mul_3486;
assign mul_4251 = slice_4249 * slice_4250;
assign slice_344 = mul_335[17:0];
assign concat_5007 = {addW_5005,slice_5006};
assign subW_1100 = subW_1099 - mul_1093;
assign slice_5763 = addW_5759[17:0];
assign lsl_1856 = add_1855 << 8;
assign slice_6519 = slice_6518[63:32];
assign add_2612 = mulnw_2609 + mulnw_2611;
assign slice_7275 = addW_7274[33:18];
assign subW_3368 = concat_3367 - concat_2815;
assign slice_4124 = slice_4123[32:16];
assign addW_217 = slice_128 + slice_30;
assign concat_4880 = {addW_4878,slice_4879};
assign subW_973 = subW_972 - mul_966;
assign slice_5636 = slice_5615[16:8];
assign mulnw_1729 = slice_1728 * slice_1725;
assign addW_6392 = slice_6387 + slice_6384;
assign mulnw_2485 = slice_2478 * slice_2484;
assign mul_7148 = slice_7146 * slice_7147;
assign lsl_3241 = add_3240 << 8;
assign slice_3997 = slice_3996[31:18];
assign slice_90 = slice_83[15:8];
assign slice_4753 = addW_4752[129:65];
assign addW_846 = slice_841 + slice_838;
assign subW_5509 = concat_5508 - concat_5448;
assign lsl_1602 = mulnw_1601 << 16;
assign addW_6265 = slice_6260 + slice_6257;
assign add_2358 = mulnw_2355 + mulnw_2357;
assign slice_7021 = slice_7020[32:16];
assign mulnw_3114 = slice_3113 * slice_3110;
assign addW_3870 = concat_3864 + subW_3869;
assign lsl_4626 = mulnw_4625 << 16;
assign add_719 = mulnw_716 + mulnw_718;
assign slice_5382 = concat_5381[63:32];
assign addW_1475 = slice_1470 + slice_1467;
assign slice_6138 = addW_6137[33:18];
assign mul_2231 = addW_2229 * addW_2230;
assign concat_6894 = {addW_6892,slice_6893};
assign concat_2987 = {addW_2985,slice_2986};
assign addW_3743 = concat_3737 + subW_3742;
assign concat_4499 = {mul_4494,slice_4498};
assign slice_592 = slice_577[7:0];
assign slice_5255 = slice_5237[15:8];
assign slice_1348 = mul_1317[15:0];
assign slice_6011 = slice_6010[31:18];
assign subW_2104 = subW_2103 - mul_2097;
assign add_6767 = lsl_6758 + add_6766;
assign addW_2860 = slice_2840 + slice_2822;
assign mul_7523 = slice_7520 * slice_7522;
assign slice_3616 = addW_3611[17:0];
assign slice_4372 = concat_4371[127:64];
assign lsl_465 = add_464 << 8;
assign slice_5128 = mul_5127[35:18];
assign slice_1221 = slice_1134[63:0];
assign subW_5884 = concat_5883 - concat_5823;
assign concat_1977 = {addW_1975,slice_1976};
assign mul_6640 = slice_6634 * slice_6636;
assign slice_2733 = slice_2727[15:0];
assign mul_7396 = slice_7392 * slice_7395;
assign mul_3489 = slice_3487 * slice_3488;
assign slice_4245 = slice_4244[31:18];
assign addW_338 = slice_333 + slice_329;
assign mul_5001 = slice_4995 * slice_4997;
assign slice_1094 = mul_1093[35:18];
assign addW_5757 = slice_5737 + slice_5696;
assign lsl_1850 = mulnw_1849 << 16;
assign subW_6513 = concat_6512 - concat_6474;
assign mulnw_2606 = slice_2604 * slice_2605;
assign concat_7269 = {addW_7267,slice_7268};
assign concat_3362 = {addW_3360,slice_3361};
assign addW_4118 = concat_4090 + addW_4117;
assign concat_211 = {concat_124,slice_210};
assign mul_4874 = slice_4868 * slice_4870;
assign slice_967 = mul_966[35:18];
assign add_5630 = mulnw_5627 + mulnw_5629;
assign add_1723 = lsl_1714 + add_1722;
assign slice_6386 = slice_6381[17:0];
assign slice_2479 = slice_2474[15:8];
assign slice_7142 = addW_7141[32:16];
assign lsl_3235 = mulnw_3234 << 16;
assign concat_3991 = {addW_3989,slice_3990};
assign mul_84 = slice_82 * slice_83;
assign addW_4747 = concat_4659 + subW_4746;
assign slice_840 = addW_835[17:0];
assign add_5503 = lsl_5501 + mul_5502;
assign mul_1596 = slice_1590 * slice_1592;
assign slice_6259 = slice_6253[17:0];
assign mulnw_2352 = slice_2350 * slice_2351;
assign slice_7015 = slice_7014[128:64];
assign add_3108 = lsl_3099 + add_3107;
assign concat_3864 = {mul_3859,slice_3863};
assign mul_4620 = slice_4618 * slice_4619;
assign mulnw_713 = slice_711 * slice_712;
assign mul_5376 = addW_5374 * addW_5375;
assign slice_1469 = addW_1464[17:0];
assign addW_6132 = concat_6126 + subW_6131;
assign slice_2225 = addW_2221[17:0];
assign mul_6888 = slice_6882 * slice_6884;
assign slice_2981 = mul_2950[15:0];
assign concat_3737 = {mul_3732,slice_3736};
assign slice_4493 = slice_4492[31:18];
assign slice_586 = mul_585[31:16];
assign mulnw_5249 = slice_5242 * slice_5248;
assign lsl_1342 = add_1341 << 8;
assign addW_6005 = concat_5999 + subW_6004;
assign slice_2098 = mul_2097[35:18];
assign slice_6761 = slice_6735[7:0];
assign slice_2854 = mul_2845[17:0];
assign slice_7517 = mul_7486[15:0];
assign concat_3610 = {concat_3590,slice_3609};
assign concat_4366 = {addW_4364,slice_4365};
assign lsl_459 = mulnw_458 << 16;
assign addW_5122 = slice_5102 + slice_5062;
assign concat_1215 = {addW_1213,slice_1214};
assign mul_5878 = addW_5876 * addW_5877;
assign slice_1971 = mul_1962[17:0];
assign slice_6634 = slice_6612[7:0];
assign slice_2727 = addW_2726[64:32];
assign slice_7390 = addW_7303[64:0];
assign slice_3483 = slice_3482[31:18];
assign add_4239 = lsl_4230 + add_4238;
assign mul_332 = slice_329 * slice_331;
assign slice_4995 = slice_4973[7:0];
assign slice_1088 = addW_1047[31:0];
assign subW_5751 = subW_5750 - mul_5744;
assign mul_1844 = slice_1838 * slice_1840;
assign mul_6507 = addW_6505 * addW_6506;
assign slice_2600 = addW_2596[15:0];
assign mul_7263 = slice_7257 * slice_7259;
assign slice_3356 = mul_3347[17:0];
assign add_4112 = mulnw_4109 + mulnw_4111;
assign subW_205 = concat_204 - concat_144;
assign slice_4868 = slice_4846[7:0];
assign slice_961 = slice_960[63:32];
assign mulnw_5624 = slice_5622 * slice_5623;
assign slice_1717 = slice_1707[7:0];
assign concat_6380 = {addW_6378,slice_6379};
assign slice_2473 = slice_2468[15:0];
assign addW_7136 = concat_7130 + subW_7135;
assign mul_3229 = slice_3223 * slice_3225;
assign slice_3985 = mul_3976[17:0];
assign addW_78 = slice_54 + slice_31;
assign subW_4741 = subW_4740 - concat_4719;
assign mulnw_5497 = slice_5496 * slice_5493;
assign slice_1590 = slice_1576[7:0];
assign slice_6253 = slice_6252[63:32];
assign slice_2346 = slice_2342[15:0];
assign subW_7009 = concat_7008 - concat_6814;
assign slice_3102 = slice_3092[7:0];
assign slice_3858 = slice_3857[31:18];
assign slice_4614 = addW_4613[32:16];
assign slice_707 = addW_703[15:0];
assign slice_5370 = slice_5366[17:0];
assign concat_1463 = {concat_1443,slice_1462};
assign concat_6126 = {mul_6121,slice_6125};
assign addW_2219 = slice_2199 + slice_2158;
assign slice_6882 = slice_6860[7:0];
assign lsl_2975 = add_2974 << 8;
assign slice_3731 = slice_3730[31:18];
assign slice_4487 = slice_4486[127:64];
assign slice_580 = slice_579[64:32];
assign slice_5243 = slice_5238[15:8];
assign lsl_1336 = mulnw_1335 << 16;
assign concat_5999 = {mul_5994,slice_5998};
assign slice_2092 = slice_2073[31:0];
assign slice_6755 = slice_6737[15:8];
assign addW_2848 = slice_2843 + slice_2839;
assign lsl_7511 = add_7510 << 8;
assign subW_3604 = mul_3603 - mul_3595;
assign mul_4360 = slice_4354 * slice_4356;
assign mul_453 = slice_447 * slice_449;
assign slice_5116 = mul_5107[17:0];
assign mul_1209 = slice_1203 * slice_1205;
assign slice_5872 = addW_5868[17:0];
assign addW_1965 = slice_1960 + slice_1956;
assign add_6628 = lsl_6626 + mul_6627;
assign addW_2721 = concat_2678 + subW_2720;
assign concat_7384 = {addW_7382,slice_7383};
assign subW_3477 = mul_3476 - mul_3468;
assign slice_4233 = slice_4207[7:0];
assign slice_326 = mul_317[17:0];
assign add_4989 = lsl_4987 + mul_4988;
assign addW_1082 = add_1068 + add_1081;
assign slice_5745 = mul_5744[35:18];
assign slice_1838 = slice_1825[7:0];
assign slice_6501 = addW_6497[17:0];
assign addW_2594 = slice_2574 + slice_2552;
assign slice_7257 = slice_7235[7:0];
assign addW_3350 = slice_3345 + slice_3341;
assign mulnw_4106 = slice_4104 * slice_4105;
assign add_199 = lsl_197 + mul_198;
assign add_4862 = lsl_4860 + mul_4861;
assign slice_955 = concat_909[31:0];
assign slice_5618 = slice_5614[15:0];
assign slice_1711 = slice_1699[16:8];
assign mul_6374 = slice_6368 * slice_6370;
assign concat_2467 = {addW_2465,slice_2466};
assign concat_7130 = {mul_7125,slice_7129};
assign slice_3223 = slice_3210[7:0];
assign addW_3979 = slice_3974 + slice_3970;
assign subW_4735 = mul_4734 - mul_4726;
assign addW_828 = add_814 + add_827;
assign add_5491 = lsl_5482 + add_5490;
assign slice_1584 = mul_1583[31:16];
assign subW_6247 = concat_6246 - concat_6186;
assign slice_2340 = slice_2339[32:16];
assign concat_7003 = {addW_7001,slice_7002};
assign slice_3096 = slice_3085[16:8];
assign addW_3852 = concat_3824 + addW_3851;
assign addW_4608 = concat_4602 + subW_4607;
assign addW_701 = slice_681 + slice_662;
assign slice_5364 = slice_5343[31:0];
assign subW_1457 = mul_1456 - mul_1448;
assign slice_6120 = slice_6119[31:18];
assign subW_2213 = subW_2212 - mul_2206;
assign add_6876 = lsl_6874 + mul_6875;
assign lsl_2969 = mulnw_2968 << 16;
assign concat_3725 = {addW_3723,slice_3724};
assign subW_4481 = concat_4480 - concat_4286;
assign addW_574 = slice_306 + slice_16;
assign slice_5237 = slice_5231[15:0];
assign mul_1330 = slice_1324 * slice_1326;
assign slice_5993 = slice_5992[31:18];
assign subW_2086 = subW_2085 - mul_2079;
assign mulnw_6749 = slice_6742 * slice_6748;
assign mul_2842 = slice_2839 * slice_2841;
assign lsl_7505 = mulnw_7504 << 16;
assign mul_3598 = slice_3596 * slice_3597;
assign slice_4354 = slice_4332[7:0];
assign slice_447 = slice_434[7:0];
assign addW_5110 = slice_5105 + slice_5101;
assign slice_1203 = slice_1181[7:0];
assign addW_5866 = slice_5824 + slice_5783;
assign mul_1959 = slice_1956 * slice_1958;
assign mulnw_6622 = slice_6621 * slice_6618;
assign addW_2715 = add_2701 + add_2714;
assign addW_7378 = slice_7373 + slice_7370;
assign mul_3471 = slice_3469 * slice_3470;
assign slice_4227 = slice_4209[15:8];
assign addW_320 = slice_315 + slice_309;
assign mulnw_4983 = slice_4982 * slice_4979;
assign mulnw_1076 = slice_1069 * slice_1075;
assign slice_5739 = slice_5698[31:0];
assign slice_1832 = mul_1831[31:16];
assign addW_6495 = slice_6475 + slice_6433;
assign subW_2588 = subW_2587 - mul_2581;
assign add_7251 = lsl_7249 + mul_7250;
assign mul_3344 = slice_3341 * slice_3343;
assign lsl_4100 = add_4099 << 8;
assign mulnw_193 = slice_192 * slice_189;
assign mulnw_4856 = slice_4855 * slice_4852;
assign addW_949 = concat_921 + addW_948;
assign addW_5612 = slice_5346 + slice_5060;
assign mul_1705 = slice_1699 * slice_1704;
assign slice_6368 = slice_6346[7:0];
assign mul_2461 = slice_2455 * slice_2457;
assign slice_7124 = slice_7123[31:18];
assign slice_3217 = mul_3216[31:16];
assign mul_3973 = slice_3970 * slice_3972;
assign subW_66 = subW_65 - mul_59;
assign mul_4729 = slice_4727 * slice_4728;
assign mulnw_822 = slice_815 * slice_821;
assign slice_5485 = slice_5475[7:0];
assign slice_1578 = addW_1577[65:33];
assign add_6241 = lsl_6239 + mul_6240;
assign subW_2334 = subW_2333 - concat_2312;
assign addW_6997 = slice_6992 + slice_6989;
assign mul_3090 = slice_3085 * slice_3089;
assign add_3846 = mulnw_3843 + mulnw_3845;
assign concat_4602 = {mul_4597,slice_4601};
assign subW_695 = subW_694 - mul_688;
assign mul_5358 = addW_5356 * addW_5357;
assign mul_1451 = slice_1449 * slice_1450;
assign addW_6114 = concat_6086 + addW_6113;
assign slice_2207 = mul_2206[35:18];
assign mulnw_6870 = slice_6869 * slice_6866;
assign mul_2963 = slice_2957 * slice_2959;
assign slice_3719 = mul_3688[15:0];
assign concat_4475 = {addW_4473,slice_4474};
assign slice_568 = concat_477[63:0];
assign slice_5231 = addW_5230[65:33];
assign slice_1324 = slice_1310[7:0];
assign concat_5987 = {addW_5985,slice_5986};
assign slice_2080 = mul_2079[35:18];
assign slice_6743 = slice_6738[15:8];
assign slice_2836 = mul_2827[17:0];
assign mul_7499 = slice_7493 * slice_7495;
assign slice_3592 = slice_3591[31:18];
assign add_4348 = lsl_4346 + mul_4347;
assign slice_441 = mul_440[31:16];
assign mul_5104 = slice_5101 * slice_5103;
assign add_1197 = lsl_1195 + mul_1196;
assign addW_5860 = add_5846 + add_5859;
assign slice_1953 = concat_1952[65:33];
assign concat_6616 = {mul_6611,slice_6615};
assign mulnw_2709 = slice_2702 * slice_2708;
assign slice_7372 = addW_7367[17:0];
assign slice_3465 = slice_3379[63:0];
assign mulnw_4221 = slice_4214 * slice_4220;
assign mul_314 = slice_309 * slice_313;
assign concat_4977 = {mul_4972,slice_4976};
assign slice_1070 = slice_1049[16:8];
assign addW_5733 = add_5719 + add_5732;
assign addW_1826 = slice_1806 + slice_1788;
assign subW_6489 = subW_6488 - mul_6482;
assign slice_2582 = mul_2581[35:18];
assign mulnw_7245 = slice_7244 * slice_7241;
assign slice_3338 = concat_3337[65:33];
assign lsl_4094 = mulnw_4093 << 16;
assign add_187 = lsl_178 + add_186;
assign concat_4850 = {mul_4845,slice_4849};
assign add_943 = mulnw_940 + mulnw_942;
assign slice_5606 = concat_5605[255:128];
assign slice_1699 = slice_1698[32:16];
assign add_6362 = lsl_6360 + mul_6361;
assign slice_2455 = slice_2433[7:0];
assign addW_7118 = concat_7112 + subW_7117;
assign addW_3211 = slice_3191 + slice_3173;
assign slice_3967 = concat_3966[63:32];
assign slice_60 = mul_59[35:18];
assign slice_4723 = addW_4722[33:18];
assign slice_816 = slice_795[16:8];
assign slice_5479 = slice_5470[16:8];
assign slice_1572 = concat_1571[127:64];
assign mulnw_6235 = slice_6234 * slice_6231;
assign subW_2328 = mul_2327 - mul_2319;
assign slice_6991 = addW_6986[17:0];
assign slice_3084 = slice_3083[64:32];
assign mulnw_3840 = slice_3838 * slice_3839;
assign slice_4596 = slice_4595[31:18];
assign slice_689 = mul_688[35:18];
assign slice_5352 = slice_5348[17:0];
assign slice_1445 = slice_1444[31:18];
assign add_6108 = mulnw_6105 + mulnw_6107;
assign slice_2201 = addW_2160[31:0];
assign concat_6864 = {mul_6859,slice_6863};
assign slice_2957 = slice_2944[7:0];
assign lsl_3713 = add_3712 << 8;
assign addW_4469 = slice_4464 + slice_4461;
assign addW_562 = concat_541 + subW_561;
assign addW_5225 = concat_5182 + subW_5224;
assign slice_1318 = mul_1317[31:16];
assign slice_5981 = mul_5950[15:0];
assign slice_2074 = slice_2073[63:32];
assign slice_6737 = slice_6729[15:0];
assign addW_2830 = slice_2825 + slice_2819;
assign slice_7493 = slice_7479[7:0];
assign add_3586 = lsl_3577 + add_3585;
assign mulnw_4342 = slice_4341 * slice_4338;
assign addW_435 = slice_415 + slice_397;
assign slice_5098 = mul_5067[15:0];
assign mulnw_1191 = slice_1190 * slice_1187;
assign mulnw_5854 = slice_5847 * slice_5853;
assign add_1947 = lsl_1945 + mul_1946;
assign slice_6610 = slice_6609[32:16];
assign slice_2703 = slice_2682[16:8];
assign concat_7366 = {concat_7346,slice_7365};
assign addW_3459 = concat_3416 + subW_3458;
assign slice_4215 = slice_4210[15:8];
assign slice_308 = slice_307[63:32];
assign slice_4971 = slice_4970[32:16];
assign add_1064 = mulnw_1061 + mulnw_1063;
assign mulnw_5727 = slice_5720 * slice_5726;
assign slice_1820 = mul_1811[17:0];
assign slice_6483 = mul_6482[35:18];
assign slice_2576 = slice_2557[31:0];
assign concat_7239 = {mul_7234,slice_7238};
assign add_3332 = lsl_3330 + mul_3331;
assign mul_4088 = slice_4086 * slice_4087;
assign slice_181 = slice_171[7:0];
assign slice_4844 = slice_4843[32:16];
assign mulnw_937 = slice_935 * slice_936;
assign concat_5600 = {addW_5598,slice_5599};
assign mulnw_6356 = slice_6355 * slice_6352;
assign add_2449 = lsl_2447 + mul_2448;
assign concat_7112 = {mul_7107,slice_7111};
assign slice_3205 = mul_3196[17:0];
assign mul_3961 = addW_3959 * addW_3960;
assign slice_54 = slice_30[31:0];
assign addW_4717 = concat_4711 + subW_4716;
assign add_810 = mulnw_807 + mulnw_809;
assign mul_5473 = slice_5470 * slice_5472;
assign concat_1566 = {addW_1564,slice_1565};
assign add_6229 = lsl_6220 + add_6228;
assign mul_2322 = slice_2320 * slice_2321;
assign concat_6985 = {concat_6943,slice_6984};
assign slice_3078 = concat_2987[63:0];
assign lsl_3834 = add_3833 << 8;
assign addW_4590 = concat_4584 + subW_4589;
assign slice_683 = slice_664[31:0];
assign slice_5346 = slice_5059[127:0];
assign add_1439 = lsl_1430 + add_1438;
assign mulnw_6102 = slice_6100 * slice_6101;
assign addW_2195 = add_2181 + add_2194;
assign slice_6858 = addW_6857[32:16];
assign slice_2951 = mul_2950[31:16];
assign lsl_3707 = mulnw_3706 << 16;
assign slice_4463 = addW_4458[17:0];
assign subW_556 = subW_555 - mul_549;
assign addW_5219 = add_5205 + add_5218;
assign slice_1312 = addW_1311[64:32];
assign lsl_5975 = add_5974 << 8;
assign slice_2068 = concat_2022[31:0];
assign addW_6731 = slice_5904 + slice_5059;
assign mul_2824 = slice_2819 * slice_2823;
assign slice_7487 = mul_7486[31:16];
assign slice_3580 = slice_3554[7:0];
assign concat_4336 = {mul_4331,slice_4335};
assign slice_429 = mul_420[17:0];
assign lsl_5092 = add_5091 << 8;
assign concat_1185 = {mul_1180,slice_1184};
assign slice_5848 = slice_5827[16:8];
assign mulnw_1941 = slice_1940 * slice_1937;
assign concat_6604 = {concat_6517,slice_6603};
assign add_2697 = mulnw_2694 + mulnw_2696;
assign subW_7360 = mul_7359 - mul_7351;
assign addW_3453 = add_3439 + add_3452;
assign slice_4209 = slice_4201[15:0];
assign subW_302 = subW_301 - concat_209;
assign addW_4965 = concat_4937 + addW_4964;
assign mulnw_1058 = slice_1056 * slice_1057;
assign slice_5721 = slice_5700[16:8];
assign addW_1814 = slice_1809 + slice_1805;
assign slice_6477 = slice_6436[31:0];
assign subW_2570 = subW_2569 - mul_2563;
assign slice_7233 = slice_7232[32:16];
assign mulnw_3326 = slice_3325 * slice_3322;
assign addW_4082 = slice_3995 + slice_3910;
assign slice_175 = slice_166[16:8];
assign concat_4838 = {addW_4836,slice_4837};
assign lsl_931 = add_930 << 8;
assign slice_5594 = mul_5585[17:0];
assign subW_1687 = subW_1686 - concat_1397;
assign concat_6350 = {mul_6345,slice_6349};
assign mulnw_2443 = slice_2442 * slice_2439;
assign slice_7106 = slice_7105[31:18];
assign addW_3199 = slice_3194 + slice_3190;
assign slice_3955 = slice_3951[17:0];
assign subW_48 = subW_47 - mul_38;
assign concat_4711 = {mul_4706,slice_4710};
assign mulnw_804 = slice_802 * slice_803;
assign slice_5467 = concat_5466[63:32];
assign mul_1560 = slice_1554 * slice_1556;
assign slice_6223 = slice_6213[7:0];
assign slice_2316 = addW_2315[33:18];
assign add_6979 = lsl_6970 + add_6978;
assign addW_3072 = concat_3051 + subW_3071;
assign lsl_3828 = mulnw_3827 << 16;
assign concat_4584 = {mul_4579,slice_4583};
assign subW_677 = subW_676 - mul_670;
assign slice_5340 = concat_5227[63:0];
assign slice_1433 = slice_1407[7:0];
assign lsl_6096 = add_6095 << 8;
assign mulnw_2189 = slice_2182 * slice_2188;
assign concat_6852 = {addW_6850,slice_6851};
assign addW_2945 = slice_2925 + slice_2907;
assign mul_3701 = slice_3695 * slice_3697;
assign concat_4457 = {concat_4415,slice_4456};
assign slice_550 = mul_549[35:18];
assign mulnw_5213 = slice_5206 * slice_5212;
assign slice_1306 = concat_1305[127:64];
assign lsl_5969 = mulnw_5968 << 16;
assign addW_2062 = concat_2034 + addW_2061;
assign slice_2818 = slice_2817[63:32];
assign slice_7481 = addW_7480[65:33];
assign slice_3574 = slice_3556[15:8];
assign slice_4330 = addW_4329[32:16];
assign addW_423 = slice_418 + slice_414;
assign lsl_5086 = mulnw_5085 << 16;
assign slice_1179 = addW_1178[32:16];
assign add_5842 = mulnw_5839 + mulnw_5841;
assign add_1935 = lsl_1926 + add_1934;
assign subW_6598 = concat_6597 - concat_6537;
assign mulnw_2691 = slice_2689 * slice_2690;
assign mul_7354 = slice_7352 * slice_7353;
assign mulnw_3447 = slice_3440 * slice_3446;
assign addW_4203 = slice_3378 + slice_2555;
assign subW_296 = concat_295 - concat_255;
assign add_4959 = mulnw_4956 + mulnw_4958;
assign slice_1052 = slice_1048[15:0];
assign add_5715 = mulnw_5712 + mulnw_5714;
assign mul_1808 = slice_1805 * slice_1807;
assign addW_6471 = add_6457 + add_6470;
assign slice_2564 = mul_2563[35:18];
assign addW_7227 = concat_7199 + addW_7226;
assign add_3320 = lsl_3311 + add_3319;
assign concat_4076 = {addW_4074,slice_4075};
assign mul_169 = slice_166 * slice_168;
assign slice_4832 = mul_4823[17:0];
assign lsl_925 = mulnw_924 << 16;
assign addW_5588 = slice_5583 + slice_5579;
assign subW_1681 = concat_1680 - concat_1486;
assign slice_6344 = slice_6343[32:16];
assign concat_2437 = {mul_2432,slice_2436};
assign concat_7100 = {addW_7098,slice_7099};
assign mul_3193 = slice_3190 * slice_3192;
assign slice_3949 = slice_3906[31:0];
assign slice_4705 = slice_4704[31:18];
assign slice_798 = slice_794[15:0];
assign mul_5461 = addW_5459 * addW_5460;
assign slice_1554 = slice_1532[7:0];
assign slice_6217 = slice_6208[16:8];
assign addW_2310 = concat_2304 + subW_2309;
assign slice_6973 = slice_6947[7:0];
assign subW_3066 = subW_3065 - mul_3059;
assign mul_3822 = slice_3820 * slice_3821;
assign slice_4578 = slice_4577[31:18];
assign slice_671 = mul_670[35:18];
assign addW_5334 = concat_5313 + subW_5333;
assign slice_1427 = slice_1409[15:8];
assign lsl_6090 = mulnw_6089 << 16;
assign slice_2183 = slice_2162[16:8];
assign addW_6846 = slice_6841 + slice_6838;
assign slice_2939 = mul_2930[17:0];
assign slice_7602 = concat_5047[511:0];
assign slice_3695 = slice_3682[7:0];
assign add_4451 = lsl_4442 + add_4450;
assign addW_544 = slice_524 + slice_484;
assign slice_5207 = slice_5186[16:8];
assign concat_1300 = {addW_1298,slice_1299};
assign mul_5963 = slice_5957 * slice_5959;
assign add_2056 = mulnw_2053 + mulnw_2055;
assign addW_6719 = concat_6430 + subW_6718;
assign subW_2812 = subW_2811 - concat_2723;
assign slice_7475 = concat_7474[129:65];
assign mulnw_3568 = slice_3561 * slice_3567;
assign concat_4324 = {addW_4322,slice_4323};
assign mul_417 = slice_414 * slice_416;
assign mul_5080 = slice_5074 * slice_5076;
assign concat_1173 = {addW_1171,slice_1172};
assign mulnw_5836 = slice_5834 * slice_5835;
assign slice_1929 = slice_1919[7:0];
assign add_6592 = lsl_6590 + mul_6591;
assign slice_2685 = addW_2681[15:0];
assign slice_7348 = slice_7347[31:18];
assign slice_3441 = slice_3420[16:8];
assign concat_4197 = {concat_3372,slice_4196};
assign mul_290 = addW_288 * addW_289;
assign mulnw_4953 = slice_4951 * slice_4952;
assign slice_1046 = slice_1045[32:16];
assign mulnw_5709 = slice_5707 * slice_5708;
assign slice_1802 = mul_1793[17:0];
assign mulnw_6465 = slice_6458 * slice_6464;
assign slice_2558 = slice_2557[63:32];
assign add_7221 = mulnw_7218 + mulnw_7220;
assign slice_3314 = slice_3304[7:0];
assign slice_4070 = mul_4039[15:0];
assign slice_163 = concat_162[63:32];
assign addW_4826 = slice_4821 + slice_4817;
assign mul_919 = slice_917 * slice_918;
assign mul_5582 = slice_5579 * slice_5581;
assign concat_1675 = {addW_1673,slice_1674};
assign concat_6338 = {concat_6251,slice_6337};
assign slice_2431 = slice_2430[32:16];
assign slice_7094 = mul_7085[17:0];
assign slice_3187 = mul_3178[17:0];
assign add_3943 = lsl_3941 + mul_3942;
assign slice_36 = slice_22[17:0];
assign addW_4699 = concat_4671 + addW_4698;
assign slice_792 = addW_750[32:0];
assign slice_5455 = slice_5451[17:0];
assign add_1548 = lsl_1546 + mul_1547;
assign mul_6211 = slice_6208 * slice_6210;
assign concat_2304 = {mul_2299,slice_2303};
assign slice_6967 = slice_6949[15:8];
assign slice_3060 = mul_3059[35:18];
assign addW_3816 = slice_3729 + slice_3644;
assign concat_4572 = {addW_4570,slice_4571};
assign slice_665 = slice_664[63:32];
assign subW_5328 = subW_5327 - mul_5321;
assign mulnw_1421 = slice_1414 * slice_1420;
assign mul_6084 = slice_6082 * slice_6083;
assign add_2177 = mulnw_2174 + mulnw_2176;
assign slice_6840 = slice_6835[17:0];
assign addW_2933 = slice_2928 + slice_2924;
assign addW_7596 = concat_6723 + subW_7595;
assign slice_3689 = mul_3688[31:16];
assign slice_4445 = slice_4419[7:0];
assign slice_538 = mul_529[17:0];
assign add_5201 = mulnw_5198 + mulnw_5200;
assign mul_1294 = slice_1288 * slice_1290;
assign slice_5957 = slice_5944[7:0];
assign mulnw_2050 = slice_2048 * slice_2049;
assign subW_6713 = subW_6712 - concat_6602;
assign subW_2806 = concat_2805 - concat_2767;
assign concat_7469 = {addW_7467,slice_7468};
assign slice_3562 = slice_3557[15:8];
assign addW_4318 = slice_4313 + slice_4310;
assign slice_411 = mul_402[17:0];
assign slice_5074 = slice_5057[7:0];
assign addW_1167 = slice_1162 + slice_1159;
assign slice_5830 = slice_5826[15:0];
assign slice_1923 = slice_1914[16:8];
assign mulnw_6586 = slice_6585 * slice_6582;
assign addW_2679 = slice_2659 + slice_2640;
assign add_7342 = lsl_7333 + add_7341;
assign add_3435 = mulnw_3432 + mulnw_3434;
assign subW_4191 = concat_4190 - concat_3638;
assign slice_284 = addW_280[17:0];
assign lsl_4947 = add_4946 << 8;
assign slice_1040 = concat_994[31:0];
assign slice_5703 = slice_5699[15:0];
assign addW_1796 = slice_1791 + slice_1786;
assign slice_6459 = slice_6438[16:8];
assign slice_2552 = slice_2551[63:32];
assign mulnw_7215 = slice_7213 * slice_7214;
assign slice_3308 = slice_3299[16:8];
assign lsl_4064 = add_4063 << 8;
assign mul_157 = addW_155 * addW_156;
assign mul_4820 = slice_4817 * slice_4819;
assign slice_913 = addW_912[32:16];
assign slice_5576 = concat_5575[63:32];
assign addW_1669 = slice_1664 + slice_1661;
assign subW_6332 = concat_6331 - concat_6271;
assign addW_7088 = slice_7083 + slice_7079;
assign addW_3181 = slice_3176 + slice_3171;
assign mulnw_3937 = slice_3936 * slice_3933;
assign slice_30 = slice_29[127:64];
assign add_4693 = mulnw_4690 + mulnw_4692;
assign add_786 = lsl_784 + mul_785;
assign slice_5449 = slice_5429[31:0];
assign mulnw_1542 = slice_1541 * slice_1538;
assign slice_6205 = concat_6204[63:32];
assign slice_2298 = slice_2297[31:18];
assign mulnw_6961 = slice_6954 * slice_6960;
assign addW_3054 = slice_3034 + slice_2994;
assign concat_3810 = {addW_3808,slice_3809};
assign slice_4566 = mul_4535[15:0];
assign slice_659 = concat_635[31:0];
assign slice_5322 = mul_5321[35:18];
assign slice_1415 = slice_1410[15:8];
assign addW_6078 = slice_5991 + slice_5906;
assign mulnw_2171 = slice_2169 * slice_2170;
assign concat_6834 = {addW_6832,slice_6833};
assign mul_2927 = slice_2924 * slice_2926;
assign subW_7590 = subW_7589 - concat_7299;
assign addW_3683 = slice_3663 + slice_3645;
assign slice_4439 = slice_4421[15:8];
assign addW_532 = slice_527 + slice_523;
assign mulnw_5195 = slice_5193 * slice_5194;
assign slice_1288 = slice_1266[7:0];
assign slice_5951 = mul_5950[31:16];
assign lsl_2044 = add_2043 << 8;
assign subW_6707 = concat_6706 - concat_6646;
assign mul_2800 = addW_2798 * addW_2799;
assign addW_7463 = slice_7458 + slice_7455;
assign slice_3556 = slice_3550[15:0];
assign slice_4312 = slice_4307[17:0];
assign addW_405 = slice_400 + slice_395;
assign slice_5068 = mul_5067[31:16];
assign slice_1161 = slice_1156[17:0];
assign slice_5824 = addW_5782[32:0];
assign mul_1917 = slice_1914 * slice_1916;
assign add_6580 = lsl_6571 + add_6579;
assign subW_2673 = subW_2672 - mul_2666;
assign slice_7336 = slice_7310[7:0];
assign mulnw_3429 = slice_3427 * slice_3428;
assign concat_4185 = {addW_4183,slice_4184};
assign addW_278 = slice_256 + slice_215;
assign lsl_4941 = mulnw_4940 << 16;
assign addW_1034 = concat_1006 + addW_1033;
assign slice_5697 = slice_5696[32:16];
assign mul_1790 = slice_1786 * slice_1789;
assign add_6453 = mulnw_6450 + mulnw_6452;
assign slice_2546 = concat_1690[255:0];
assign lsl_7209 = add_7208 << 8;
assign mul_3302 = slice_3299 * slice_3301;
assign lsl_4058 = mulnw_4057 << 16;
assign slice_151 = slice_147[17:0];
assign slice_4814 = concat_4813[63:32];
assign addW_907 = concat_901 + subW_906;
assign mul_5570 = addW_5568 * addW_5569;
assign slice_1663 = addW_1658[17:0];
assign add_6326 = lsl_6324 + mul_6325;
assign subW_2419 = subW_2418 - concat_2397;
assign mul_7082 = slice_7079 * slice_7081;
assign mul_3175 = slice_3171 * slice_3174;
assign add_3931 = lsl_3922 + add_3930;
assign mulnw_4687 = slice_4685 * slice_4686;
assign mulnw_780 = slice_779 * slice_776;
assign mul_5443 = addW_5441 * addW_5442;
assign concat_1536 = {mul_1531,slice_1535};
assign mul_6199 = addW_6197 * addW_6198;
assign addW_2292 = concat_2264 + addW_2291;
assign slice_6955 = slice_6950[15:8];
assign slice_3048 = mul_3039[17:0];
assign slice_3804 = mul_3773[15:0];
assign lsl_4560 = add_4559 << 8;
assign addW_653 = concat_647 + subW_652;
assign addW_5316 = slice_5274 + slice_5234;
assign slice_1409 = slice_1402[15:0];
assign concat_6072 = {addW_6070,slice_6071};
assign slice_2165 = slice_2161[15:0];
assign addW_6828 = slice_6823 + slice_6820;
assign slice_2921 = mul_2912[17:0];
assign subW_7584 = concat_7583 - concat_7389;
assign slice_3677 = mul_3668[17:0];
assign mulnw_4433 = slice_4426 * slice_4432;
assign mul_526 = slice_523 * slice_525;
assign slice_5189 = addW_5185[15:0];
assign add_1282 = lsl_1280 + mul_1281;
assign addW_5945 = slice_5925 + slice_5907;
assign lsl_2038 = mulnw_2037 << 16;
assign mul_6701 = addW_6699 * addW_6700;
assign slice_2794 = addW_2790[17:0];
assign slice_7457 = addW_7452[17:0];
assign slice_3550 = addW_3549[64:32];
assign concat_4306 = {addW_4304,slice_4305};
assign mul_399 = slice_395 * slice_398;
assign slice_5062 = slice_5061[64:32];
assign concat_1155 = {addW_1153,slice_1154};
assign add_5818 = lsl_5816 + mul_5817;
assign slice_1911 = mul_1880[15:0];
assign slice_6574 = slice_6564[7:0];
assign slice_2667 = mul_2666[35:18];
assign slice_7330 = slice_7312[15:8];
assign slice_3423 = addW_3419[15:0];
assign slice_4179 = mul_4170[17:0];
assign slice_272 = mul_263[17:0];
assign mul_4935 = slice_4933 * slice_4934;
assign add_1028 = mulnw_1025 + mulnw_1027;
assign subW_5691 = subW_5690 - concat_5669;
assign slice_1784 = slice_1696[63:0];
assign mulnw_6447 = slice_6445 * slice_6446;
assign addW_2540 = concat_2248 + subW_2539;
assign lsl_7203 = mulnw_7202 << 16;
assign slice_3296 = mul_3265[15:0];
assign mul_4052 = slice_4046 * slice_4048;
assign slice_145 = slice_125[31:0];
assign mul_4808 = addW_4806 * addW_4807;
assign concat_901 = {mul_896,slice_900};
assign slice_5564 = slice_5560[17:0];
assign concat_1657 = {concat_1615,slice_1656};
assign mulnw_6320 = slice_6319 * slice_6316;
assign subW_2413 = mul_2412 - mul_2404;
assign slice_7076 = concat_7075[63:32];
assign slice_3169 = addW_3082[63:0];
assign slice_3925 = slice_3915[7:0];
assign lsl_4681 = add_4680 << 8;
assign add_774 = lsl_765 + add_773;
assign slice_5437 = slice_5433[17:0];
assign slice_1530 = addW_1529[32:16];
assign slice_6193 = slice_6189[17:0];
assign add_2286 = mulnw_2283 + mulnw_2285;
assign slice_6949 = slice_6944[15:0];
assign addW_3042 = slice_3037 + slice_3033;
assign lsl_3798 = add_3797 << 8;
assign lsl_4554 = mulnw_4553 << 16;
assign concat_647 = {mul_642,slice_646};
assign slice_5310 = mul_5279[15:0];
assign slice_1403 = slice_1402[32:16];
assign slice_6066 = mul_6035[15:0];
assign slice_2159 = slice_2158[32:16];
assign slice_6822 = slice_6816[17:0];
assign addW_2915 = slice_2910 + slice_2905;
assign concat_7578 = {addW_7576,slice_7577};
assign addW_3671 = slice_3666 + slice_3662;
assign slice_4427 = slice_4422[15:8];
assign slice_520 = mul_489[15:0];
assign addW_5183 = slice_5163 + slice_5144;
assign mulnw_1276 = slice_1275 * slice_1272;
assign slice_5939 = mul_5930[17:0];
assign mul_2032 = slice_2030 * slice_2031;
assign slice_6695 = addW_6691[17:0];
assign addW_2788 = slice_2768 + slice_2727;
assign concat_7451 = {concat_7431,slice_7450};
assign addW_3544 = concat_3501 + subW_3543;
assign addW_4300 = slice_4295 + slice_4292;
assign slice_393 = slice_306[63:0];
assign slice_5056 = slice_5055[64:32];
assign addW_1149 = slice_1144 + slice_1141;
assign mulnw_5812 = slice_5811 * slice_5808;
assign lsl_1905 = add_1904 << 8;
assign slice_6568 = slice_6559[16:8];
assign slice_2661 = slice_2642[31:0];
assign mulnw_7324 = slice_7317 * slice_7323;
assign addW_3417 = slice_3397 + slice_3376;
assign addW_4173 = slice_4168 + slice_4164;
assign addW_266 = slice_261 + slice_257;
assign addW_4929 = slice_4842 + slice_4757;
assign mulnw_1022 = slice_1020 * slice_1021;
assign subW_5685 = mul_5684 - mul_5676;
assign concat_1778 = {addW_1776,slice_1777};
assign slice_6441 = slice_6437[15:0];
assign subW_2534 = subW_2533 - concat_2422;
assign mul_7197 = slice_7195 * slice_7196;
assign lsl_3290 = add_3289 << 8;
assign slice_4046 = slice_4033[7:0];
assign mul_139 = addW_137 * addW_138;
assign slice_4802 = slice_4798[17:0];
assign slice_895 = slice_894[31:18];
assign slice_5558 = addW_5516[31:0];
assign add_1651 = lsl_1642 + add_1650;
assign add_6314 = lsl_6305 + add_6313;
assign mul_2407 = slice_2405 * slice_2406;
assign mul_7070 = addW_7068 * addW_7069;
assign concat_3163 = {addW_3161,slice_3162};
assign slice_3919 = slice_3908[16:8];
assign lsl_4675 = mulnw_4674 << 16;
assign slice_768 = slice_758[7:0];
assign slice_5431 = slice_5430[31:18];
assign concat_1524 = {addW_1522,slice_1523};
assign slice_6187 = slice_6166[31:0];
assign mulnw_2280 = slice_2278 * slice_2279;
assign concat_6943 = {addW_6941,slice_6942};
assign mul_3036 = slice_3033 * slice_3035;
assign lsl_3792 = mulnw_3791 << 16;
assign mul_4548 = slice_4542 * slice_4544;
assign slice_641 = addW_640[33:18];
assign lsl_5304 = add_5303 << 8;
assign concat_1397 = {addW_1395,slice_1396};
assign lsl_6060 = add_6059 << 8;
assign slice_2153 = concat_2107[31:0];
assign slice_6816 = slice_6815[63:32];
assign mul_2909 = slice_2905 * slice_2908;
assign addW_7572 = slice_7567 + slice_7564;
assign mul_3665 = slice_3662 * slice_3664;
assign slice_4421 = slice_4416[15:0];
assign lsl_514 = add_513 << 8;
assign subW_5177 = subW_5176 - mul_5170;
assign concat_1270 = {mul_1265,slice_1269};
assign addW_5933 = slice_5928 + slice_5924;
assign slice_2026 = addW_2025[32:16];
assign addW_6689 = slice_6647 + slice_6606;
assign subW_2782 = subW_2781 - mul_2775;
assign subW_7445 = mul_7444 - mul_7436;
assign addW_3538 = add_3524 + add_3537;
assign slice_4294 = slice_4288[17:0];
assign concat_387 = {addW_385,slice_386};
assign slice_1143 = slice_1136[17:0];
assign add_5806 = lsl_5797 + add_5805;
assign lsl_1899 = mulnw_1898 << 16;
assign mul_6562 = slice_6559 * slice_6561;
assign subW_2655 = subW_2654 - mul_2648;
assign slice_7318 = slice_7313[15:8];
assign subW_3411 = subW_3410 - mul_3404;
assign mul_4167 = slice_4164 * slice_4166;
assign mul_260 = slice_257 * slice_259;
assign concat_4923 = {addW_4921,slice_4922};
assign lsl_1016 = add_1015 << 8;
assign mul_5679 = slice_5677 * slice_5678;
assign addW_1772 = slice_1767 + slice_1764;
assign addW_6435 = slice_6169 + slice_5905;
assign subW_2528 = concat_2527 - concat_2467;
assign addW_7191 = slice_7104 + slice_7019;
assign lsl_3284 = mulnw_3283 << 16;
assign slice_4040 = mul_4039[31:16];
assign slice_133 = slice_129[17:0];
assign slice_4796 = slice_4753[31:0];
assign addW_889 = concat_883 + subW_888;
assign add_5552 = lsl_5550 + mul_5551;
assign slice_1645 = slice_1619[7:0];
assign slice_6308 = slice_6298[7:0];
assign slice_2401 = addW_2400[33:18];
assign slice_7064 = slice_7060[17:0];
assign addW_3157 = slice_3152 + slice_3149;
assign mul_3913 = slice_3908 * slice_3912;
assign mul_4669 = slice_4667 * slice_4668;
assign slice_762 = slice_752[16:8];
assign subW_5425 = subW_5424 - concat_5381;
assign addW_1518 = slice_1513 + slice_1510;
assign mul_6181 = addW_6179 * addW_6180;
assign lsl_2274 = add_2273 << 8;
assign mul_6937 = slice_6931 * slice_6933;
assign slice_3030 = mul_2999[15:0];
assign mul_3786 = slice_3780 * slice_3782;
assign slice_4542 = slice_4529[7:0];
assign concat_635 = {addW_633,slice_634};
assign lsl_5298 = mulnw_5297 << 16;
assign slice_1391 = concat_1367[31:0];
assign lsl_6054 = mulnw_6053 << 16;
assign addW_2147 = concat_2119 + addW_2146;
assign subW_6810 = concat_6809 - concat_6771;
assign slice_2903 = slice_2816[63:0];
assign slice_7566 = addW_7561[17:0];
assign slice_3659 = mul_3650[17:0];
assign concat_4415 = {addW_4413,slice_4414};
assign lsl_508 = mulnw_507 << 16;
assign slice_5171 = mul_5170[35:18];
assign slice_1264 = addW_1263[32:16];
assign mul_5927 = slice_5924 * slice_5926;
assign addW_2020 = concat_2014 + subW_2019;
assign addW_6683 = add_6669 + add_6682;
assign slice_2776 = mul_2775[35:18];
assign mul_7439 = slice_7437 * slice_7438;
assign mulnw_3532 = slice_3525 * slice_3531;
assign slice_4288 = slice_4287[63:32];
assign mul_381 = slice_375 * slice_377;
assign subW_5044 = subW_5043 - concat_4195;
assign slice_1137 = slice_1136[31:18];
assign slice_5800 = slice_5790[7:0];
assign mul_1893 = slice_1887 * slice_1889;
assign slice_6556 = concat_6555[63:32];
assign slice_2649 = mul_2648[35:18];
assign slice_7312 = slice_7305[15:0];
assign slice_3405 = mul_3404[35:18];
assign slice_4161 = concat_4160[65:33];
assign slice_254 = mul_223[15:0];
assign slice_4917 = mul_4908[17:0];
assign lsl_1010 = mulnw_1009 << 16;
assign slice_5673 = addW_5672[33:18];
assign slice_1766 = addW_1761[17:0];
assign slice_6429 = concat_6428[255:128];
assign mul_2522 = addW_2520 * addW_2521;
assign concat_7185 = {addW_7183,slice_7184};
assign mul_3278 = slice_3272 * slice_3274;
assign addW_4034 = slice_4014 + slice_3996;
assign slice_127 = slice_126[31:18];
assign add_4790 = lsl_4788 + mul_4789;
assign concat_883 = {mul_878,slice_882};
assign mulnw_5546 = slice_5545 * slice_5542;
assign slice_1639 = slice_1621[15:8];
assign slice_6302 = slice_6293[16:8];
assign addW_2395 = concat_2389 + subW_2394;
assign slice_7058 = slice_7015[31:0];
assign slice_3151 = addW_3146[17:0];
assign slice_3907 = slice_3906[64:32];
assign OUTPUT = concat_7603;
    endmodule